**************************************************
* Manufacturer:          Würth Elektronik
* Kinds:                 MLCCs Capacitors
* Matchcode:             WCAP-CSGP
* Library Type:          LTspice
* Version:               rev22c
* Created/modified by:   Ella
* Date and Time:         10/13/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 0402_885012105004_470nF 1 2
Rser 1 3 0.0135620044546
Lser 2 4 2.89834924E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0402_885012105004_470nF
*******
.subckt 0402_885012105005_680nF 1 2
Rser 1 3 0.00866869355558
Lser 2 4 3.2312296E-10
C1 3 4 0.00000068
Rpar 3 4 200000000
.ends 0402_885012105005_680nF
*******
.subckt 0402_885012105006_1uF 1 2
Rser 1 3 0.0122136788791
Lser 2 4 3.38680925E-10
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0402_885012105006_1uF
*******
.subckt 0402_885012105007_2.2uF 1 2
Rser 1 3 0.00909909650012
Lser 2 4 3.49876612E-10
C1 3 4 0.0000022
Rpar 3 4 20000000
.ends 0402_885012105007_2.2uF
*******
.subckt 0402_885012105008_4.7uF 1 2
Rser 1 3 0.00453732146966
Lser 2 4 3.78498478E-10
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0402_885012105008_4.7uF
*******
.subckt 0402_885012105020_10uF 1 2
Rser 1 3 0.0058
Lser 2 4 0.0000000008
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0402_885012105020_10uF
*******
.subckt 0603_885012106001_470nF 1 2
Rser 1 3 0.00946787785536
Lser 2 4 2.50326617E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0603_885012106001_470nF
*******
.subckt 0603_885012106002_680nF 1 2
Rser 1 3 0.0104592893966
Lser 2 4 3.4734058E-10
C1 3 4 0.00000068
Rpar 3 4 200000000
.ends 0603_885012106002_680nF
*******
.subckt 0603_885012106003_1uF 1 2
Rser 1 3 0.00760558670624
Lser 2 4 3.54495768E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012106003_1uF
*******
.subckt 0603_885012106004_2.2uF 1 2
Rser 1 3 0.00652337052819
Lser 2 4 4.58001637E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0603_885012106004_2.2uF
*******
.subckt 0603_885012106005_4.7uF 1 2
Rser 1 3 0.00436564105168
Lser 2 4 5.20484374E-10
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0603_885012106005_4.7uF
*******
.subckt 0603_885012106006_10uF 1 2
Rser 1 3 0.00407641026021
Lser 2 4 4.16060333E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0603_885012106006_10uF
*******
.subckt 0805_885012107001_2.2uF 1 2
Rser 1 3 0.00487002224398
Lser 2 4 2.50543345E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012107001_2.2uF
*******
.subckt 0805_885012107002_3.3uF 1 2
Rser 1 3 0.00453837206006
Lser 2 4 2.98091685E-10
C1 3 4 0.0000033
Rpar 3 4 30000000
.ends 0805_885012107002_3.3uF
*******
.subckt 0805_885012107003_4.7uF 1 2
Rser 1 3 0.00422571742874
Lser 2 4 2.56201535E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0805_885012107003_4.7uF
*******
.subckt 0805_885012107004_10uF 1 2
Rser 1 3 0.00320609856405
Lser 2 4 3.83098838E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 0805_885012107004_10uF
*******
.subckt 0805_885012107005_22uF 1 2
Rser 1 3 0.00282261758127
Lser 2 4 5.44199046E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 0805_885012107005_22uF
*******
.subckt 0805_885012107006_47uF 1 2
Rser 1 3 0.00246814753418
Lser 2 4 4.62831333E-10
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 0805_885012107006_47uF
*******
.subckt 1206_885012108001_4.7uF 1 2
Rser 1 3 0.00600320174513
Lser 2 4 5.14564007E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012108001_4.7uF
*******
.subckt 1206_885012108002_10uF 1 2
Rser 1 3 0.00340980665018
Lser 2 4 8.40328091E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012108002_10uF
*******
.subckt 1206_885012108003_22uF 1 2
Rser 1 3 0.003095358264
Lser 2 4 8.67209117E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1206_885012108003_22uF
*******
.subckt 1206_885012108004_47uF 1 2
Rser 1 3 0.00304958303174
Lser 2 4 8.27626832E-10
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1206_885012108004_47uF
*******
.subckt 1206_885012108005_100uF 1 2
Rser 1 3 0.00189819698397
Lser 2 4 0.0000000009
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 1206_885012108005_100uF
*******
.subckt 1210_885012109001_10uF 1 2
Rser 1 3 0.00236975905543
Lser 2 4 7.97405226E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1210_885012109001_10uF
*******
.subckt 1210_885012109002_22uF 1 2
Rser 1 3 0.00298875292394
Lser 2 4 0.0000000009
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1210_885012109002_22uF
*******
.subckt 1210_885012109003_47uF 1 2
Rser 1 3 0.00230591969867
Lser 2 4 9.5617691E-10
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1210_885012109003_47uF
*******
.subckt 1210_885012109004_100uF 1 2
Rser 1 3 0.00239801642091
Lser 2 4 0.0000000009
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 1210_885012109004_100uF
*******
.subckt 0603_885012206001_470nF 1 2
Rser 1 3 0.00945
Lser 2 4 0.00000000041822
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0603_885012206001_470nF
*******
.subckt 0603_885012206002_1uF 1 2
Rser 1 3 0.00781
Lser 2 4 0.00000000043943
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012206002_1uF
*******
.subckt 0805_885012207001_2.2uF 1 2
Rser 1 3 0.00442275214815
Lser 2 4 2.37717125E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012207001_2.2uF
*******
.subckt 0805_885012207002_4.7uF 1 2
Rser 1 3 0.00447387150505
Lser 2 4 2.50863578E-10
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0805_885012207002_4.7uF
*******
.subckt 0805_885012207003_10uF 1 2
Rser 1 3 0.00336648172245
Lser 2 4 4.89291579E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0805_885012207003_10uF
*******
.subckt 1206_885012208001_2.2uF 1 2
Rser 1 3 0.00708971442636
Lser 2 4 4.50708422E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 1206_885012208001_2.2uF
*******
.subckt 1206_885012208002_4.7uF 1 2
Rser 1 3 0.00380516684832
Lser 2 4 4.86025433E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012208002_4.7uF
*******
.subckt 1206_885012208003_10uF 1 2
Rser 1 3 0.00257769589302
Lser 2 4 7.50158848E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012208003_10uF
*******
.subckt 0201_885012104003_100nF 1 2
Rser 1 3 0.02829
Lser 2 4 0.00000000018
C1 3 4 0.0000001
Rpar 3 4 500000000
.ends 0201_885012104003_100nF
*******
.subckt 0201_885012104004_10nF 1 2
Rser 1 3 0.0627
Lser 2 4 0.000000000218
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012104004_10nF
*******
.subckt 0201_885012104009_100nF 1 2
Rser 1 3 0.0337
Lser 2 4 0.00000000018
C1 3 4 0.0000001
Rpar 3 4 500000000
.ends 0201_885012104009_100nF
*******
.subckt 0201_885012104010_220nF 1 2
Rser 1 3 0.043
Lser 2 4 0.00000000021
C1 3 4 0.00000022
Rpar 3 4 200000000
.ends 0201_885012104010_220nF
*******
.subckt 0201_885012104011_1uF 1 2
Rser 1 3 0.0109
Lser 2 4 0.00000000023
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0201_885012104011_1uF
*******
.subckt 0402_885012005049_1pF 1 2
Rser 1 3 0.372412566115
Lser 2 4 3.42487064E-10
C1 3 4 0.000000000001
Rpar 3 4 10000000000
.ends 0402_885012005049_1pF
*******
.subckt 0402_885012005050_1.5pF 1 2
Rser 1 3 0.262794296584
Lser 2 4 3.57764917E-10
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0402_885012005050_1.5pF
*******
.subckt 0402_885012005051_2.2pF 1 2
Rser 1 3 0.373107051593
Lser 2 4 3.52926651E-10
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0402_885012005051_2.2pF
*******
.subckt 0402_885012005052_3.3pF 1 2
Rser 1 3 0.371592714575
Lser 2 4 3.85528579E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0402_885012005052_3.3pF
*******
.subckt 0402_885012005053_4.7pF 1 2
Rser 1 3 0.443688812845
Lser 2 4 4.55408482E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0402_885012005053_4.7pF
*******
.subckt 0402_885012005054_6.8pF 1 2
Rser 1 3 0.397780736645
Lser 2 4 4.18761945E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0402_885012005054_6.8pF
*******
.subckt 0402_885012005055_10pF 1 2
Rser 1 3 0.367986500147
Lser 2 4 4.54592782E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005055_10pF
*******
.subckt 0402_885012005056_15pF 1 2
Rser 1 3 0.289002377009
Lser 2 4 4.35524241E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885012005056_15pF
*******
.subckt 0402_885012005057_22pF 1 2
Rser 1 3 0.1946461244
Lser 2 4 4.43759844E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885012005057_22pF
*******
.subckt 0402_885012005058_33pF 1 2
Rser 1 3 0.125165063018
Lser 2 4 4.11479308E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005058_33pF
*******
.subckt 0402_885012005059_47pF 1 2
Rser 1 3 0.136483462277
Lser 2 4 4.44322285E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005059_47pF
*******
.subckt 0402_885012005060_68pF 1 2
Rser 1 3 0.101411214779
Lser 2 4 4.24748886E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005060_68pF
*******
.subckt 0402_885012005061_100pF 1 2
Rser 1 3 0.0708016190464
Lser 2 4 3.72654022E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005061_100pF
*******
.subckt 0402_885012005062_150pF 1 2
Rser 1 3 0.043551770519
Lser 2 4 3.72165147E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012005062_150pF
*******
.subckt 0402_885012005063_220pF 1 2
Rser 1 3 0.0328677075671
Lser 2 4 3.55619232E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012005063_220pF
*******
.subckt 0402_885012005067_1nF 1 2
Rser 1 3 0.065
Lser 2 4 0.000000001
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012005067_1nF
*******
.subckt 0603_885012006048_3.3pF 1 2
Rser 1 3 0.351777802818
Lser 2 4 4.93521689E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0603_885012006048_3.3pF
*******
.subckt 0603_885012006049_4.7pF 1 2
Rser 1 3 0.314951809581
Lser 2 4 4.34213899E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0603_885012006049_4.7pF
*******
.subckt 0603_885012006050_6.8pF 1 2
Rser 1 3 0.53
Lser 2 4 0.00000000049
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0603_885012006050_6.8pF
*******
.subckt 0603_885012006051_10pF 1 2
Rser 1 3 0.423568844547
Lser 2 4 6.08699424E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006051_10pF
*******
.subckt 0603_885012006052_15pF 1 2
Rser 1 3 0.396040749585
Lser 2 4 6.08298711E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006052_15pF
*******
.subckt 0603_885012006053_22pF 1 2
Rser 1 3 0.388744823765
Lser 2 4 6.9588017E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006053_22pF
*******
.subckt 0603_885012006054_33pF 1 2
Rser 1 3 0.321193198235
Lser 2 4 7.31689517E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006054_33pF
*******
.subckt 0603_885012006055_47pF 1 2
Rser 1 3 0.290935011258
Lser 2 4 4.02698987E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006055_47pF
*******
.subckt 0603_885012006056_68pF 1 2
Rser 1 3 0.190199312239
Lser 2 4 6.75111985E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006056_68pF
*******
.subckt 0603_885012006057_100pF 1 2
Rser 1 3 0.155626039874
Lser 2 4 4.37579661E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006057_100pF
*******
.subckt 0603_885012006058_150pF 1 2
Rser 1 3 0.117171082106
Lser 2 4 5.86950362E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006058_150pF
*******
.subckt 0603_885012006059_220pF 1 2
Rser 1 3 0.120673949599
Lser 2 4 6.11171216E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012006059_220pF
*******
.subckt 0603_885012006060_330pF 1 2
Rser 1 3 0.0984499950001
Lser 2 4 5.75039775E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006060_330pF
*******
.subckt 0603_885012006061_470pF 1 2
Rser 1 3 0.0701665420081
Lser 2 4 5.55279727E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006061_470pF
*******
.subckt 0603_885012006062_680pF 1 2
Rser 1 3 0.058780576404
Lser 2 4 5.07120306E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006062_680pF
*******
.subckt 0603_885012006063_1nF 1 2
Rser 1 3 0.040317449025
Lser 2 4 4.45418718E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006063_1nF
*******
.subckt 0805_885012007046_1.5pF 1 2
Rser 1 3 0.498754904967
Lser 2 4 4.46307458E-10
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0805_885012007046_1.5pF
*******
.subckt 0805_885012007047_2.2pF 1 2
Rser 1 3 0.464027184378
Lser 2 4 4.17958974E-10
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0805_885012007047_2.2pF
*******
.subckt 0805_885012007048_3.3pF 1 2
Rser 1 3 0.476983731701
Lser 2 4 4.57833988E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0805_885012007048_3.3pF
*******
.subckt 0805_885012007049_4.7pF 1 2
Rser 1 3 0.497100489266
Lser 2 4 4.97943432E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0805_885012007049_4.7pF
*******
.subckt 0805_885012007050_6.8pF 1 2
Rser 1 3 0.437292047874
Lser 2 4 5.43803179E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0805_885012007050_6.8pF
*******
.subckt 0805_885012007051_10pF 1 2
Rser 1 3 0.5317
Lser 2 4 0.00000000045
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0805_885012007051_10pF
*******
.subckt 0805_885012007052_15pF 1 2
Rser 1 3 0.351715326777
Lser 2 4 5.44262413E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007052_15pF
*******
.subckt 0805_885012007053_22pF 1 2
Rser 1 3 0.320807516938
Lser 2 4 5.98353392E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0805_885012007053_22pF
*******
.subckt 0805_885012007054_33pF 1 2
Rser 1 3 0.251170142371
Lser 2 4 5.67157711E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007054_33pF
*******
.subckt 0805_885012007055_47pF 1 2
Rser 1 3 0.216515950035
Lser 2 4 5.20835554E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885012007055_47pF
*******
.subckt 0805_885012007056_68pF 1 2
Rser 1 3 0.173987704202
Lser 2 4 4.36318354E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0805_885012007056_68pF
*******
.subckt 0805_885012007057_100pF 1 2
Rser 1 3 0.112239658687
Lser 2 4 3.23857063E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007057_100pF
*******
.subckt 0805_885012007058_150pF 1 2
Rser 1 3 0.125944924272
Lser 2 4 4.46129224E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007058_150pF
*******
.subckt 0805_885012007059_220pF 1 2
Rser 1 3 0.079249932999
Lser 2 4 3.92377309E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012007059_220pF
*******
.subckt 0805_885012007060_330pF 1 2
Rser 1 3 0.0873115639161
Lser 2 4 4.48869509E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007060_330pF
*******
.subckt 0805_885012007061_470pF 1 2
Rser 1 3 0.0447460793708
Lser 2 4 5.13925095E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007061_470pF
*******
.subckt 0805_885012007062_680pF 1 2
Rser 1 3 0.0641329981739
Lser 2 4 4.25300517E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012007062_680pF
*******
.subckt 0805_885012007063_1nF 1 2
Rser 1 3 0.0594421507531
Lser 2 4 4.12205624E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007063_1nF
*******
.subckt 0805_885012007064_1.5nF 1 2
Rser 1 3 0.0542761813318
Lser 2 4 4.44523189E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012007064_1.5nF
*******
.subckt 0805_885012007065_2.2nF 1 2
Rser 1 3 0.0452125293188
Lser 2 4 3.18286842E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012007065_2.2nF
*******
.subckt 0805_885012007066_3.3nF 1 2
Rser 1 3 0.0386718470366
Lser 2 4 4.52637868E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012007066_3.3nF
*******
.subckt 0805_885012007067_4.7nF 1 2
Rser 1 3 0.0321239026517
Lser 2 4 3.90170133E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012007067_4.7nF
*******
.subckt 1206_885012008037_10pF 1 2
Rser 1 3 0.247786722229
Lser 2 4 5.75498755E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1206_885012008037_10pF
*******
.subckt 1206_885012008038_15pF 1 2
Rser 1 3 0.203981995296
Lser 2 4 5.79093876E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 1206_885012008038_15pF
*******
.subckt 1206_885012008039_22pF 1 2
Rser 1 3 0.160102464353
Lser 2 4 5.19970978E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1206_885012008039_22pF
*******
.subckt 1206_885012008040_33pF 1 2
Rser 1 3 0.211299340525
Lser 2 4 5.80360065E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 1206_885012008040_33pF
*******
.subckt 1206_885012008041_47pF 1 2
Rser 1 3 0.208069659743
Lser 2 4 5.31192815E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885012008041_47pF
*******
.subckt 1206_885012008042_68pF 1 2
Rser 1 3 0.207112222887
Lser 2 4 5.32291452E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 1206_885012008042_68pF
*******
.subckt 1206_885012008043_100pF 1 2
Rser 1 3 0.120593750684
Lser 2 4 4.75662979E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008043_100pF
*******
.subckt 1206_885012008044_150pF 1 2
Rser 1 3 0.116934479556
Lser 2 4 4.79036564E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012008044_150pF
*******
.subckt 1206_885012008045_220pF 1 2
Rser 1 3 0.10386657318
Lser 2 4 4.26569823E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012008045_220pF
*******
.subckt 1206_885012008046_330pF 1 2
Rser 1 3 0.0889473100116
Lser 2 4 3.86799658E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012008046_330pF
*******
.subckt 1206_885012008047_470pF 1 2
Rser 1 3 0.112293156509
Lser 2 4 4.49592146E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012008047_470pF
*******
.subckt 1206_885012008048_680pF 1 2
Rser 1 3 0.0885483556492
Lser 2 4 4.83404689E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012008048_680pF
*******
.subckt 1206_885012008049_1nF 1 2
Rser 1 3 0.0678258865879
Lser 2 4 4.38251746E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012008049_1nF
*******
.subckt 1206_885012008050_1.5nF 1 2
Rser 1 3 0.0522994987595
Lser 2 4 3.90875574E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012008050_1.5nF
*******
.subckt 1206_885012008051_2.2nF 1 2
Rser 1 3 0.0481287677862
Lser 2 4 4.23334149E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012008051_2.2nF
*******
.subckt 1206_885012008052_3.3nF 1 2
Rser 1 3 0.048551433153
Lser 2 4 3.89367659E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012008052_3.3nF
*******
.subckt 1206_885012008053_4.7nF 1 2
Rser 1 3 0.0373751695173
Lser 2 4 3.96656883E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012008053_4.7nF
*******
.subckt 1206_885012008054_6.8nF 1 2
Rser 1 3 0.0328755784645
Lser 2 4 4.18880071E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008054_6.8nF
*******
.subckt 1206_885012008055_10nF 1 2
Rser 1 3 0.0308699044735
Lser 2 4 4.5821325E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008055_10nF
*******
.subckt 1210_885012009007_22pF 1 2
Rser 1 3 0.374121714519
Lser 2 4 2.35270135E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1210_885012009007_22pF
*******
.subckt 1210_885012009008_33pF 1 2
Rser 1 3 0.242364797292
Lser 2 4 2.04183536E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 1210_885012009008_33pF
*******
.subckt 1210_885012009009_47pF 1 2
Rser 1 3 0.210290362797
Lser 2 4 2.1842961E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1210_885012009009_47pF
*******
.subckt 1210_885012009010_68pF 1 2
Rser 1 3 0.147762447298
Lser 2 4 1.90656729E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 1210_885012009010_68pF
*******
.subckt 1210_885012009011_100pF 1 2
Rser 1 3 0.129347366442
Lser 2 4 2.02608781E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1210_885012009011_100pF
*******
.subckt 1210_885012009012_150pF 1 2
Rser 1 3 0.130052835884
Lser 2 4 2.16784494E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1210_885012009012_150pF
*******
.subckt 1210_885012009013_220pF 1 2
Rser 1 3 0.0421105658392
Lser 2 4 2.03486371E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1210_885012009013_220pF
*******
.subckt 1210_885012009014_330pF 1 2
Rser 1 3 0.0366680474844
Lser 2 4 2.12935248E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1210_885012009014_330pF
*******
.subckt 1210_885012009015_470pF 1 2
Rser 1 3 0.041753756573
Lser 2 4 3.51053092E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1210_885012009015_470pF
*******
.subckt 1210_885012009016_680pF 1 2
Rser 1 3 0.0310627645209
Lser 2 4 2.06977272E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1210_885012009016_680pF
*******
.subckt 1210_885012009017_1nF 1 2
Rser 1 3 0.0212060307253
Lser 2 4 2.0371621E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885012009017_1nF
*******
.subckt 1210_885012009018_1.5nF 1 2
Rser 1 3 0.0312392079081
Lser 2 4 2.87207915E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1210_885012009018_1.5nF
*******
.subckt 1210_885012009019_2.2nF 1 2
Rser 1 3 0.0215418747712
Lser 2 4 2.06777607E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1210_885012009019_2.2nF
*******
.subckt 1210_885012009020_3.3nF 1 2
Rser 1 3 0.0267047192368
Lser 2 4 2.05676794E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1210_885012009020_3.3nF
*******
.subckt 1210_885012009021_4.7nF 1 2
Rser 1 3 0.0311921178887
Lser 2 4 2.6092549E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1210_885012009021_4.7nF
*******
.subckt 1210_885012009022_6.8nF 1 2
Rser 1 3 0.0328474651911
Lser 2 4 1.68986675E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1210_885012009022_6.8nF
*******
.subckt 1210_885012009023_10nF 1 2
Rser 1 3 0.0123831418384
Lser 2 4 1.88456734E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1210_885012009023_10nF
*******
.subckt 1210_885012009024_15nF 1 2
Rser 1 3 0.0151582048451
Lser 2 4 2.71190675E-10
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1210_885012009024_15nF
*******
.subckt 1812_885012010005_100pF 1 2
Rser 1 3 0.12355169432
Lser 2 4 3.51203653E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1812_885012010005_100pF
*******
.subckt 1812_885012010006_220pF 1 2
Rser 1 3 0.0878558292315
Lser 2 4 3.98601571E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1812_885012010006_220pF
*******
.subckt 1812_885012010007_470pF 1 2
Rser 1 3 0.0486179980779
Lser 2 4 3.42708418E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1812_885012010007_470pF
*******
.subckt 1812_885012010008_1nF 1 2
Rser 1 3 0.054974361057
Lser 2 4 3.20553197E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_885012010008_1nF
*******
.subckt 1812_885012010009_1.5nF 1 2
Rser 1 3 0.0235411944876
Lser 2 4 3.17035352E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1812_885012010009_1.5nF
*******
.subckt 1812_885012010010_3.3nF 1 2
Rser 1 3 0.0199944630408
Lser 2 4 3.02916593E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1812_885012010010_3.3nF
*******
.subckt 1812_885012010011_4.7nF 1 2
Rser 1 3 0.0944854934425
Lser 2 4 4.17148603E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1812_885012010011_4.7nF
*******
.subckt 1812_885012010012_6.8nF 1 2
Rser 1 3 0.0862794087323
Lser 2 4 2.93234437E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1812_885012010012_6.8nF
*******
.subckt 1812_885012010013_10nF 1 2
Rser 1 3 0.0378661246646
Lser 2 4 3.63058436E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012010013_10nF
*******
.subckt 1812_885012010014_15nF 1 2
Rser 1 3 0.0258373805332
Lser 2 4 2.604228E-10
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1812_885012010014_15nF
*******
.subckt 1812_885012010015_22nF 1 2
Rser 1 3 0.0255141881395
Lser 2 4 3.80015608E-10
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1812_885012010015_22nF
*******
.subckt 1812_885012010016_33nF 1 2
Rser 1 3 0.0536968994705
Lser 2 4 3.37435968E-10
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1812_885012010016_33nF
*******
.subckt 1206_885012108022_10uF 1 2
Rser 1 3 0.00342327531378
Lser 2 4 0.000000000799
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012108022_10uF
*******
.subckt 0402_885012205055_100pF 1 2
Rser 1 3 0.81826
Lser 2 4 0.00000000027428
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012205055_100pF
*******
.subckt 0402_885012205056_150pF 1 2
Rser 1 3 0.632711426036
Lser 2 4 1.20280732E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012205056_150pF
*******
.subckt 0402_885012205057_220pF 1 2
Rser 1 3 0.578964014005
Lser 2 4 1.69232145E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012205057_220pF
*******
.subckt 0402_885012205058_330pF 1 2
Rser 1 3 0.503553103715
Lser 2 4 1.67673778E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012205058_330pF
*******
.subckt 0402_885012205059_470pF 1 2
Rser 1 3 0.341891187733
Lser 2 4 1.53352894E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012205059_470pF
*******
.subckt 0402_885012205060_680pF 1 2
Rser 1 3 0.291776877274
Lser 2 4 1.90727531E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0402_885012205060_680pF
*******
.subckt 0402_885012205061_1nF 1 2
Rser 1 3 0.16682
Lser 2 4 0.00000000027542
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205061_1nF
*******
.subckt 0402_885012205062_1.5nF 1 2
Rser 1 3 0.318149132739
Lser 2 4 2.00030416E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0402_885012205062_1.5nF
*******
.subckt 0402_885012205063_2.2nF 1 2
Rser 1 3 0.167940534432
Lser 2 4 1.9652905E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0402_885012205063_2.2nF
*******
.subckt 0402_885012205064_3.3nF 1 2
Rser 1 3 0.128032535119
Lser 2 4 2.21229721E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0402_885012205064_3.3nF
*******
.subckt 0402_885012205065_4.7nF 1 2
Rser 1 3 0.12665496656
Lser 2 4 2.40553052E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205065_4.7nF
*******
.subckt 0402_885012205066_6.8nF 1 2
Rser 1 3 0.103789689499
Lser 2 4 1.90645336E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0402_885012205066_6.8nF
*******
.subckt 0402_885012205067_10nF 1 2
Rser 1 3 0.110942181295
Lser 2 4 1.63617133E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0402_885012205067_10nF
*******
.subckt 0402_885012205086_100nF 1 2
Rser 1 3 0.07
Lser 2 4 0.00000000055
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0402_885012205086_100nF
*******
.subckt 0402_885012205092_100nF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000006
C1 3 4 0.0000001
Rpar 3 4 500000000
.ends 0402_885012205092_100nF
*******
.subckt 0603_885012206077_100pF 1 2
Rser 1 3 0.85996
Lser 2 4 0.00000000023099
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206077_100pF
*******
.subckt 0603_885012206078_150pF 1 2
Rser 1 3 0.6711
Lser 2 4 0.00000000028059
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012206078_150pF
*******
.subckt 0603_885012206079_220pF 1 2
Rser 1 3 0.58208
Lser 2 4 0.00000000030164
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012206079_220pF
*******
.subckt 0603_885012206080_330pF 1 2
Rser 1 3 0.43473
Lser 2 4 0.00000000032084
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206080_330pF
*******
.subckt 0603_885012206081_470pF 1 2
Rser 1 3 0.34619
Lser 2 4 0.00000000032738
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206081_470pF
*******
.subckt 0603_885012206082_680pF 1 2
Rser 1 3 0.303992916785
Lser 2 4 3.80425244E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206082_680pF
*******
.subckt 0603_885012206083_1nF 1 2
Rser 1 3 0.25783718447
Lser 2 4 4.104475E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206083_1nF
*******
.subckt 0603_885012206083R_1nF 1 2
Rser 1 3 0.25783718447
Lser 2 4 4.104475E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206083R_1nF
*******
.subckt 0603_885012206084_1.5nF 1 2
Rser 1 3 0.180999474852
Lser 2 4 3.54773595E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206084_1.5nF
*******
.subckt 0603_885012206085_2.2nF 1 2
Rser 1 3 0.139424404216
Lser 2 4 3.27512531E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012206085_2.2nF
*******
.subckt 0603_885012206086_3.3nF 1 2
Rser 1 3 0.105745225203
Lser 2 4 3.39462116E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206086_3.3nF
*******
.subckt 0603_885012206087_4.7nF 1 2
Rser 1 3 0.0821607581427
Lser 2 4 2.83989011E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206087_4.7nF
*******
.subckt 0603_885012206088_6.8nF 1 2
Rser 1 3 0.0838686105847
Lser 2 4 4.16447222E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206088_6.8nF
*******
.subckt 0603_885012206089_10nF 1 2
Rser 1 3 0.0358532866879
Lser 2 4 3.4059544E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206089_10nF
*******
.subckt 0603_885012206089R_10nF 1 2
Rser 1 3 0.0358532866879
Lser 2 4 3.4059544E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206089R_10nF
*******
.subckt 0603_885012206090_15nF 1 2
Rser 1 3 0.0485012368007
Lser 2 4 3.32575255E-10
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0603_885012206090_15nF
*******
.subckt 0603_885012206091_22nF 1 2
Rser 1 3 0.00971971773084
Lser 2 4 3.00225265E-10
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885012206091_22nF
*******
.subckt 0603_885012206092_33nF 1 2
Rser 1 3 0.02322
Lser 2 4 0.00000000030071
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0603_885012206092_33nF
*******
.subckt 0603_885012206093_47nF 1 2
Rser 1 3 0.02723
Lser 2 4 0.00000000027891
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0603_885012206093_47nF
*******
.subckt 0603_885012206094_68nF 1 2
Rser 1 3 0.01852
Lser 2 4 0.00000000023609
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0603_885012206094_68nF
*******
.subckt 0603_885012206095_100nF 1 2
Rser 1 3 0.0157659152881
Lser 2 4 3.10171966E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206095_100nF
*******
.subckt 0603_885012206095R_100nF 1 2
Rser 1 3 0.0157659152881
Lser 2 4 3.10171966E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206095R_100nF
*******
.subckt 0603_885012206121_330nF 1 2
Rser 1 3 0.0116331902783
Lser 2 4 2.98906197E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012206121_330nF
*******
.subckt 0603_885012206125_220nF 1 2
Rser 1 3 0.017
Lser 2 4 0.000000001
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012206125_220nF
*******
.subckt 0805_885012207080_100pF 1 2
Rser 1 3 0.88248
Lser 2 4 0.00000000026383
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207080_100pF
*******
.subckt 0805_885012207081_150pF 1 2
Rser 1 3 0.74128
Lser 2 4 0.00000000030962
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012207081_150pF
*******
.subckt 0805_885012207082_220pF 1 2
Rser 1 3 0.48326
Lser 2 4 0.00000000027382
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012207082_220pF
*******
.subckt 0805_885012207083_330pF 1 2
Rser 1 3 0.40314
Lser 2 4 0.00000000028019
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012207083_330pF
*******
.subckt 0805_885012207084_470pF 1 2
Rser 1 3 0.29801
Lser 2 4 0.00000000032037
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207084_470pF
*******
.subckt 0805_885012207085_680pF 1 2
Rser 1 3 0.24191
Lser 2 4 0.00000000035763
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012207085_680pF
*******
.subckt 0805_885012207086_1nF 1 2
Rser 1 3 0.16468
Lser 2 4 0.00000000030011
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207086_1nF
*******
.subckt 0805_885012207087_1.5nF 1 2
Rser 1 3 0.14696
Lser 2 4 0.00000000040084
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207087_1.5nF
*******
.subckt 0805_885012207088_2.2nF 1 2
Rser 1 3 0.11179
Lser 2 4 0.00000000038067
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012207088_2.2nF
*******
.subckt 0805_885012207089_3.3nF 1 2
Rser 1 3 0.08492
Lser 2 4 0.0000000003695
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207089_3.3nF
*******
.subckt 0805_885012207090_4.7nF 1 2
Rser 1 3 0.05225
Lser 2 4 0.00000000025076
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012207090_4.7nF
*******
.subckt 0805_885012207091_6.8nF 1 2
Rser 1 3 0.06481
Lser 2 4 0.00000000034495
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0805_885012207091_6.8nF
*******
.subckt 0805_885012207092_10nF 1 2
Rser 1 3 0.06275
Lser 2 4 0.00000000031024
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207092_10nF
*******
.subckt 0805_885012207093_15nF 1 2
Rser 1 3 0.04594
Lser 2 4 0.00000000031216
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0805_885012207093_15nF
*******
.subckt 0805_885012207094_22nF 1 2
Rser 1 3 0.04966
Lser 2 4 0.00000000031956
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0805_885012207094_22nF
*******
.subckt 0805_885012207095_33nF 1 2
Rser 1 3 0.0344549798517
Lser 2 4 0.00000000043
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0805_885012207095_33nF
*******
.subckt 0805_885012207096_47nF 1 2
Rser 1 3 0.0256748827303
Lser 2 4 0.00000000038
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0805_885012207096_47nF
*******
.subckt 0805_885012207097_68nF 1 2
Rser 1 3 0.0207501013107
Lser 2 4 0.00000000038
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0805_885012207097_68nF
*******
.subckt 0805_885012207098_100nF 1 2
Rser 1 3 0.0175748078756
Lser 2 4 0.0000000004
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207098_100nF
*******
.subckt 0805_885012207098R_100nF 1 2
Rser 1 3 0.0175748078756
Lser 2 4 0.0000000004
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207098R_100nF
*******
.subckt 0805_885012207099_150nF 1 2
Rser 1 3 0.0142447362747
Lser 2 4 0.00000000045
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0805_885012207099_150nF
*******
.subckt 0805_885012207100_220nF 1 2
Rser 1 3 0.0120359560176
Lser 2 4 0.00000000044
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885012207100_220nF
*******
.subckt 0805_885012207101_330nF 1 2
Rser 1 3 0.0111899844274
Lser 2 4 0.00000000048
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885012207101_330nF
*******
.subckt 0805_885012207102_470nF 1 2
Rser 1 3 0.00874819634126
Lser 2 4 0.000000000465
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0805_885012207102_470nF
*******
.subckt 0805_885012207103_1uF 1 2
Rser 1 3 0.0053065272233
Lser 2 4 2.83466289E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0805_885012207103_1uF
*******
.subckt 0805_885012207103R_1uF 1 2
Rser 1 3 0.0053065272233
Lser 2 4 2.83466289E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0805_885012207103R_1uF
*******
.subckt 1206_885012208070_150pF 1 2
Rser 1 3 0.71274
Lser 2 4 0.00000000032053
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012208070_150pF
*******
.subckt 1206_885012208071_220pF 1 2
Rser 1 3 0.50529569726
Lser 2 4 2.96273344E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012208071_220pF
*******
.subckt 1206_885012208072_330pF 1 2
Rser 1 3 0.43202
Lser 2 4 0.00000000057877
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012208072_330pF
*******
.subckt 1206_885012208073_470pF 1 2
Rser 1 3 0.34146
Lser 2 4 0.00000000040636
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208073_470pF
*******
.subckt 1206_885012208074_680pF 1 2
Rser 1 3 0.34068
Lser 2 4 0.00000000050397
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012208074_680pF
*******
.subckt 1206_885012208075_1nF 1 2
Rser 1 3 0.22519
Lser 2 4 0.00000000041699
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208075_1nF
*******
.subckt 1206_885012208076_1.5nF 1 2
Rser 1 3 0.18074
Lser 2 4 0.00000000040041
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012208076_1.5nF
*******
.subckt 1206_885012208077_2.2nF 1 2
Rser 1 3 0.13842
Lser 2 4 0.00000000039067
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012208077_2.2nF
*******
.subckt 1206_885012208078_3.3nF 1 2
Rser 1 3 0.13733
Lser 2 4 0.00000000045693
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012208078_3.3nF
*******
.subckt 1206_885012208079_4.7nF 1 2
Rser 1 3 0.09403
Lser 2 4 0.00000000040583
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208079_4.7nF
*******
.subckt 1206_885012208080_6.8nF 1 2
Rser 1 3 0.08271
Lser 2 4 0.00000000048076
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012208080_6.8nF
*******
.subckt 1206_885012208081_10nF 1 2
Rser 1 3 0.07548
Lser 2 4 0.00000000050044
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208081_10nF
*******
.subckt 1206_885012208082_15nF 1 2
Rser 1 3 0.06346
Lser 2 4 0.00000000050869
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1206_885012208082_15nF
*******
.subckt 1206_885012208083_22nF 1 2
Rser 1 3 0.05996
Lser 2 4 0.00000000050024
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1206_885012208083_22nF
*******
.subckt 1206_885012208084_33nF 1 2
Rser 1 3 0.07214
Lser 2 4 0.00000000048096
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1206_885012208084_33nF
*******
.subckt 1206_885012208085_47nF 1 2
Rser 1 3 0.05144
Lser 2 4 0.00000000044024
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1206_885012208085_47nF
*******
.subckt 1206_885012208086_68nF 1 2
Rser 1 3 0.03887
Lser 2 4 0.00000000042372
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 1206_885012208086_68nF
*******
.subckt 1206_885012208087_100nF 1 2
Rser 1 3 0.02357
Lser 2 4 0.00000000059109
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885012208087_100nF
*******
.subckt 1206_885012208088_150nF 1 2
Rser 1 3 0.01669
Lser 2 4 0.00000000057596
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1206_885012208088_150nF
*******
.subckt 1206_885012208089_220nF 1 2
Rser 1 3 0.01154
Lser 2 4 0.0000000005471
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1206_885012208089_220nF
*******
.subckt 1206_885012208090_330nF 1 2
Rser 1 3 0.01154
Lser 2 4 0.00000000068941
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1206_885012208090_330nF
*******
.subckt 1206_885012208091_470nF 1 2
Rser 1 3 0.01065
Lser 2 4 0.00000000073215
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1206_885012208091_470nF
*******
.subckt 1206_885012208092_680nF 1 2
Rser 1 3 0.00829
Lser 2 4 0.00000000068878
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1206_885012208092_680nF
*******
.subckt 1206_885012208093_1uF 1 2
Rser 1 3 0.00556
Lser 2 4 0.00000000059996
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885012208093_1uF
*******
.subckt 1206_885012208094_4.7uF 1 2
Rser 1 3 0.00352
Lser 2 4 0.00000000057332
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012208094_4.7uF
*******
.subckt 1210_885012209029_1nF 1 2
Rser 1 3 0.24578
Lser 2 4 0.00000000010314
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885012209029_1nF
*******
.subckt 1210_885012209030_1.5nF 1 2
Rser 1 3 0.21363
Lser 2 4 0.00000000011258
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1210_885012209030_1.5nF
*******
.subckt 1210_885012209031_2.2nF 1 2
Rser 1 3 0.17328
Lser 2 4 0.00000000013551
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1210_885012209031_2.2nF
*******
.subckt 1210_885012209032_3.3nF 1 2
Rser 1 3 0.10148
Lser 2 4 0.000000000079128
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1210_885012209032_3.3nF
*******
.subckt 1210_885012209033_4.7nF 1 2
Rser 1 3 0.12905
Lser 2 4 0.00000000012069
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1210_885012209033_4.7nF
*******
.subckt 1210_885012209034_6.8nF 1 2
Rser 1 3 0.05767
Lser 2 4 0.0000000001329
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1210_885012209034_6.8nF
*******
.subckt 1210_885012209035_10nF 1 2
Rser 1 3 0.07029
Lser 2 4 0.00000000063234
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1210_885012209035_10nF
*******
.subckt 1210_885012209036_15nF 1 2
Rser 1 3 0.04823
Lser 2 4 0.00000000065476
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1210_885012209036_15nF
*******
.subckt 1210_885012209037_22nF 1 2
Rser 1 3 0.0318
Lser 2 4 0.0000000005907
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1210_885012209037_22nF
*******
.subckt 1210_885012209038_33nF 1 2
Rser 1 3 0.02862
Lser 2 4 0.00000000012573
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1210_885012209038_33nF
*******
.subckt 1210_885012209039_47nF 1 2
Rser 1 3 0.01636
Lser 2 4 0.00000000055283
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1210_885012209039_47nF
*******
.subckt 1210_885012209040_68nF 1 2
Rser 1 3 0.02967
Lser 2 4 0.00000000066933
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 1210_885012209040_68nF
*******
.subckt 1210_885012209041_100nF 1 2
Rser 1 3 0.0232640980559
Lser 2 4 5.50483551E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1210_885012209041_100nF
*******
.subckt 1210_885012209042_150nF 1 2
Rser 1 3 0.0151905172405
Lser 2 4 5.27589443E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1210_885012209042_150nF
*******
.subckt 1210_885012209043_220nF 1 2
Rser 1 3 0.0127857665848
Lser 2 4 5.1481312E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1210_885012209043_220nF
*******
.subckt 1210_885012209044_330nF 1 2
Rser 1 3 0.00839371610696
Lser 2 4 5.53587415E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1210_885012209044_330nF
*******
.subckt 1210_885012209045_470nF 1 2
Rser 1 3 0.00675106116736
Lser 2 4 5.53881923E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1210_885012209045_470nF
*******
.subckt 1210_885012209046_680nF 1 2
Rser 1 3 0.00595213609047
Lser 2 4 5.69870142E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1210_885012209046_680nF
*******
.subckt 1210_885012209047_1uF 1 2
Rser 1 3 0.0444403254894
Lser 2 4 7.99001148E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209047_1uF
*******
.subckt 1210_885012209047R_1uF 1 2
Rser 1 3 0.0444403254894
Lser 2 4 7.99001148E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209047R_1uF
*******
.subckt 1210_885012209048_4.7uF 1 2
Rser 1 3 0.00278836774782
Lser 2 4 2.60340728E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1210_885012209048_4.7uF
*******
.subckt 1210_885012209073_10uF 1 2
Rser 1 3 0.00803494307495
Lser 2 4 4.01881911E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1210_885012209073_10uF
*******
.subckt 1812_885012210013_1nF 1 2
Rser 1 3 0.22122
Lser 2 4 0.00000000021688
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_885012210013_1nF
*******
.subckt 1812_885012210014_1.5nF 1 2
Rser 1 3 0.17474
Lser 2 4 0.00000000020664
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1812_885012210014_1.5nF
*******
.subckt 1812_885012210015_2.2nF 1 2
Rser 1 3 0.13333
Lser 2 4 0.00000000015464
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1812_885012210015_2.2nF
*******
.subckt 1812_885012210016_3.3nF 1 2
Rser 1 3 0.11987
Lser 2 4 0.00000000054219
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1812_885012210016_3.3nF
*******
.subckt 1812_885012210017_4.7nF 1 2
Rser 1 3 0.08329
Lser 2 4 0.00000000014772
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1812_885012210017_4.7nF
*******
.subckt 1812_885012210018_6.8nF 1 2
Rser 1 3 0.08602
Lser 2 4 0.00000000061736
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1812_885012210018_6.8nF
*******
.subckt 1812_885012210019_10nF 1 2
Rser 1 3 0.07293
Lser 2 4 0.00000000052871
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012210019_10nF
*******
.subckt 1812_885012210020_15nF 1 2
Rser 1 3 0.067
Lser 2 4 0.0000000007302
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1812_885012210020_15nF
*******
.subckt 1812_885012210021_22nF 1 2
Rser 1 3 0.05662
Lser 2 4 0.00000000062074
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1812_885012210021_22nF
*******
.subckt 1812_885012210022_33nF 1 2
Rser 1 3 0.03888
Lser 2 4 0.00000000053993
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1812_885012210022_33nF
*******
.subckt 1812_885012210023_47nF 1 2
Rser 1 3 0.0333
Lser 2 4 0.00000000024107
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1812_885012210023_47nF
*******
.subckt 1812_885012210024_68nF 1 2
Rser 1 3 0.0283
Lser 2 4 0.00000000079079
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 1812_885012210024_68nF
*******
.subckt 1812_885012210025_100nF 1 2
Rser 1 3 0.0434286733285
Lser 2 4 5.51116314E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1812_885012210025_100nF
*******
.subckt 1812_885012210026_150nF 1 2
Rser 1 3 0.0274984909595
Lser 2 4 6.78013757E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1812_885012210026_150nF
*******
.subckt 1812_885012210027_220nF 1 2
Rser 1 3 0.0210915166325
Lser 2 4 5.00831292E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1812_885012210027_220nF
*******
.subckt 1812_885012210028_330nF 1 2
Rser 1 3 0.0146375735099
Lser 2 4 4.50409847E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1812_885012210028_330nF
*******
.subckt 1812_885012210029_470nF 1 2
Rser 1 3 0.0117735855692
Lser 2 4 3.80795098E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1812_885012210029_470nF
*******
.subckt 1812_885012210030_680nF 1 2
Rser 1 3 0.00705429391862
Lser 2 4 4.5048548E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1812_885012210030_680nF
*******
.subckt 1812_885012210031_1uF 1 2
Rser 1 3 0.00507618175382
Lser 2 4 5.00373592E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1812_885012210031_1uF
*******
.subckt 1812_885012210032_2.2uF 1 2
Rser 1 3 0.00377371050938
Lser 2 4 4.19292053E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1812_885012210032_2.2uF
*******
.subckt 0201_885012204001_100pF 1 2
Rser 1 3 0.8951
Lser 2 4 0.00000000017
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0201_885012204001_100pF
*******
.subckt 0201_885012204002_680pF 1 2
Rser 1 3 0.3189
Lser 2 4 0.00000000022
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0201_885012204002_680pF
*******
.subckt 0201_885012204003_1nF 1 2
Rser 1 3 0.2506
Lser 2 4 0.00000000021
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0201_885012204003_1nF
*******
.subckt 0201_885012004002_47pF 1 2
Rser 1 3 0.2226
Lser 2 4 0.0000000002
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0201_885012004002_47pF
*******
.subckt 0201_885012004011_10pF 1 2
Rser 1 3 0.5169
Lser 2 4 0.00000000022
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0201_885012004011_10pF
*******
.subckt 0201_885012004012_22pF 1 2
Rser 1 3 0.4505
Lser 2 4 0.000000000253
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0201_885012004012_22pF
*******
.subckt 0201_885012004013_33pF 1 2
Rser 1 3 0.2722
Lser 2 4 0.00000000022
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0201_885012004013_33pF
*******
.subckt 0201_885012004014_100pF 1 2
Rser 1 3 0.1789
Lser 2 4 0.0000000002
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0201_885012004014_100pF
*******
.subckt 2220_885012214005_10uF 1 2
Rser 1 3 0.003
Lser 2 4 0.0000000012
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 2220_885012214005_10uF
*******
.subckt 0603_885012206126_1uF 1 2
Rser 1 3 0.0115
Lser 2 4 0.0000000008
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0603_885012206126_1uF
*******
.subckt 0402_885012005074_10pF 1 2
Rser 1 3 0.421651463477
Lser 2 4 4.14790783E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005074_10pF
*******
.subckt 0402_885012005077_33pF 1 2
Rser 1 3 0.221604982314
Lser 2 4 3.49022204E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005077_33pF
*******
.subckt 0402_885012005078_47pF 1 2
Rser 1 3 0.24210526915
Lser 2 4 4.45579658E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005078_47pF
*******
.subckt 0402_885012005079_68pF 1 2
Rser 1 3 0.204212177962
Lser 2 4 3.70169713E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005079_68pF
*******
.subckt 0402_885012005080_100pF 1 2
Rser 1 3 0.117553952575
Lser 2 4 3.96667338E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005080_100pF
*******
.subckt 0402_885012005085_8.2pF 1 2
Rser 1 3 0.352598551895
Lser 2 4 4.16869039E-10
C1 3 4 0.0000000000082
Rpar 3 4 10000000000
.ends 0402_885012005085_8.2pF
*******
.subckt 0603_885012006073_10pF 1 2
Rser 1 3 0.407424144741
Lser 2 4 5.41304078E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006073_10pF
*******
.subckt 0603_885012006074_15pF 1 2
Rser 1 3 0.380584852252
Lser 2 4 5.65804545E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006074_15pF
*******
.subckt 0603_885012006076_33pF 1 2
Rser 1 3 0.286862998414
Lser 2 4 6.50561095E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006076_33pF
*******
.subckt 0603_885012006077_47pF 1 2
Rser 1 3 0.245803082005
Lser 2 4 6.35972597E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006077_47pF
*******
.subckt 0603_885012006078_68pF 1 2
Rser 1 3 0.200732636434
Lser 2 4 5.98671906E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006078_68pF
*******
.subckt 0603_885012006079_100pF 1 2
Rser 1 3 0.147736548124
Lser 2 4 5.50713639E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006079_100pF
*******
.subckt 0603_885012006080_150pF 1 2
Rser 1 3 0.123096464746
Lser 2 4 5.27226081E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006080_150pF
*******
.subckt 0603_885012006082_330pF 1 2
Rser 1 3 0.0953300210797
Lser 2 4 4.24072373E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006082_330pF
*******
.subckt 0603_885012006083_470pF 1 2
Rser 1 3 0.0701382798145
Lser 2 4 4.13398494E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006083_470pF
*******
.subckt 0603_885012006084_680pF 1 2
Rser 1 3 0.0621072894488
Lser 2 4 4.13475086E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006084_680pF
*******
.subckt 0603_885012006085_1nF 1 2
Rser 1 3 0.0532527583524
Lser 2 4 3.27557981E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006085_1nF
*******
.subckt 0805_885012007076_10pF 1 2
Rser 1 3 0.348978588999
Lser 2 4 4.65201661E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0805_885012007076_10pF
*******
.subckt 0805_885012007077_15pF 1 2
Rser 1 3 0.299948487506
Lser 2 4 4.54423504E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007077_15pF
*******
.subckt 0805_885012007079_33pF 1 2
Rser 1 3 0.121980282644
Lser 2 4 4.43859848E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007079_33pF
*******
.subckt 0805_885012007080_47pF 1 2
Rser 1 3 0.166811229395
Lser 2 4 4.10637959E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885012007080_47pF
*******
.subckt 0805_885012007081_68pF 1 2
Rser 1 3 0.180760159531
Lser 2 4 3.86267029E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0805_885012007081_68pF
*******
.subckt 0805_885012007082_100pF 1 2
Rser 1 3 0.0753079048439
Lser 2 4 2.90973988E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007082_100pF
*******
.subckt 0805_885012007083_150pF 1 2
Rser 1 3 0.198942265358
Lser 2 4 3.89898948E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007083_150pF
*******
.subckt 0805_885012007085_330pF 1 2
Rser 1 3 0.0776936134254
Lser 2 4 2.60803415E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007085_330pF
*******
.subckt 0805_885012007086_470pF 1 2
Rser 1 3 0.0588553647502
Lser 2 4 2.97840521E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007086_470pF
*******
.subckt 0805_885012007087_680pF 1 2
Rser 1 3 0.0627822674091
Lser 2 4 2.56856486E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012007087_680pF
*******
.subckt 0805_885012007088_1nF 1 2
Rser 1 3 0.0369190815603
Lser 2 4 3.02824205E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007088_1nF
*******
.subckt 0805_885012007089_1.5nF 1 2
Rser 1 3 0.0444913409463
Lser 2 4 3.70041338E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012007089_1.5nF
*******
.subckt 0805_885012007091_3.3nF 1 2
Rser 1 3 0.0238862333296
Lser 2 4 3.52340361E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012007091_3.3nF
*******
.subckt 0805_885012007092_4.7nF 1 2
Rser 1 3 0.0360290329923
Lser 2 4 3.13853583E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012007092_4.7nF
*******
.subckt 1206_885012008061_10pF 1 2
Rser 1 3 0.375598705152
Lser 2 4 5.61558997E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1206_885012008061_10pF
*******
.subckt 1206_885012008062_15pF 1 2
Rser 1 3 0.35
Lser 2 4 0.00000000056
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 1206_885012008062_15pF
*******
.subckt 1206_885012008065_47pF 1 2
Rser 1 3 0.19407783985
Lser 2 4 5.43052823E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885012008065_47pF
*******
.subckt 1206_885012008067_100pF 1 2
Rser 1 3 0.157459451422
Lser 2 4 4.64194319E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008067_100pF
*******
.subckt 1206_885012008068_150pF 1 2
Rser 1 3 0.130548247324
Lser 2 4 4.36494773E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012008068_150pF
*******
.subckt 1206_885012008070_330pF 1 2
Rser 1 3 0.0931468259828
Lser 2 4 4.33607632E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012008070_330pF
*******
.subckt 1206_885012008071_470pF 1 2
Rser 1 3 0.0863181912042
Lser 2 4 4.5763957E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012008071_470pF
*******
.subckt 1206_885012008072_680pF 1 2
Rser 1 3 0.0777497909642
Lser 2 4 4.75215911E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012008072_680pF
*******
.subckt 1206_885012008073_1nF 1 2
Rser 1 3 0.0477152917275
Lser 2 4 4.99751981E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012008073_1nF
*******
.subckt 1206_885012008074_1.5nF 1 2
Rser 1 3 0.0354598757287
Lser 2 4 3.99445906E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012008074_1.5nF
*******
.subckt 1206_885012008076_3.3nF 1 2
Rser 1 3 0.0314389546323
Lser 2 4 4.34527012E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012008076_3.3nF
*******
.subckt 1206_885012008078_6.8nF 1 2
Rser 1 3 0.0257323206072
Lser 2 4 4.35781903E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008078_6.8nF
*******
.subckt 1206_885012008079_10nF 1 2
Rser 1 3 0.0235458917441
Lser 2 4 4.56933086E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008079_10nF
*******
.subckt 0402_885012205080_1nF 1 2
Rser 1 3 0.25
Lser 2 4 0.00000000044
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205080_1nF
*******
.subckt 0402_885012205084_4.7nF 1 2
Rser 1 3 0.155
Lser 2 4 0.0000000004
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205084_4.7nF
*******
.subckt 0603_885012206102_100pF 1 2
Rser 1 3 0.903793201449
Lser 2 4 4.30927368E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206102_100pF
*******
.subckt 0603_885012206103_150pF 1 2
Rser 1 3 0.663307587764
Lser 2 4 4.01639305E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012206103_150pF
*******
.subckt 0603_885012206105_330pF 1 2
Rser 1 3 0.471881844186
Lser 2 4 4.17174312E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206105_330pF
*******
.subckt 0603_885012206106_470pF 1 2
Rser 1 3 0.3
Lser 2 4 0.000000000401
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206106_470pF
*******
.subckt 0603_885012206107_680pF 1 2
Rser 1 3 0.307694453707
Lser 2 4 4.68126223E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206107_680pF
*******
.subckt 0603_885012206108_1nF 1 2
Rser 1 3 0.202024514637
Lser 2 4 5.1469819E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206108_1nF
*******
.subckt 0603_885012206109_1.5nF 1 2
Rser 1 3 0.160907873586
Lser 2 4 4.36594994E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206109_1.5nF
*******
.subckt 0603_885012206111_3.3nF 1 2
Rser 1 3 0.141390340152
Lser 2 4 5.69446762E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206111_3.3nF
*******
.subckt 0603_885012206112_4.7nF 1 2
Rser 1 3 0.0887774662878
Lser 2 4 4.3949757E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206112_4.7nF
*******
.subckt 0603_885012206113_6.8nF 1 2
Rser 1 3 0.0566471875739
Lser 2 4 4.04270889E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206113_6.8nF
*******
.subckt 0603_885012206114_10nF 1 2
Rser 1 3 0.0614305159536
Lser 2 4 4.58570264E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206114_10nF
*******
.subckt 0603_885012206114R_10nF 1 2
Rser 1 3 0.0614305159536
Lser 2 4 4.58570264E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206114R_10nF
*******
.subckt 0603_885012206118_47nF 1 2
Rser 1 3 0.0260966431276
Lser 2 4 4.02961106E-10
C1 3 4 0.000000047
Rpar 3 4 2100000000
.ends 0603_885012206118_47nF
*******
.subckt 0603_885012206120_100nF 1 2
Rser 1 3 0.02
Lser 2 4 0.0000000008
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0603_885012206120_100nF
*******
.subckt 0805_885012207110_100pF 1 2
Rser 1 3 0.893542107954
Lser 2 4 3.72840309E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207110_100pF
*******
.subckt 0805_885012207111_150pF 1 2
Rser 1 3 0.75393192763
Lser 2 4 4.30786527E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012207111_150pF
*******
.subckt 0805_885012207113_330pF 1 2
Rser 1 3 0.884149804092
Lser 2 4 3.16830341E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012207113_330pF
*******
.subckt 0805_885012207114_470pF 1 2
Rser 1 3 0.374236748173
Lser 2 4 4.69987959E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207114_470pF
*******
.subckt 0805_885012207115_680pF 1 2
Rser 1 3 0.441399652418
Lser 2 4 3.85533833E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012207115_680pF
*******
.subckt 0805_885012207116_1nF 1 2
Rser 1 3 0.200201288389
Lser 2 4 4.27706413E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207116_1nF
*******
.subckt 0805_885012207117_1.5nF 1 2
Rser 1 3 0.165813253283
Lser 2 4 4.70069305E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207117_1.5nF
*******
.subckt 0805_885012207119_3.3nF 1 2
Rser 1 3 0.107994017051
Lser 2 4 4.67027278E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207119_3.3nF
*******
.subckt 0805_885012207120_4.7nF 1 2
Rser 1 3 0.0819387083384
Lser 2 4 4.01268553E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012207120_4.7nF
*******
.subckt 0805_885012207121_6.8nF 1 2
Rser 1 3 0.0730376666068
Lser 2 4 4.71078792E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0805_885012207121_6.8nF
*******
.subckt 0805_885012207122_10nF 1 2
Rser 1 3 0.0602542793423
Lser 2 4 5.20580851E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207122_10nF
*******
.subckt 0805_885012207123_15nF 1 2
Rser 1 3 0.0418698831686
Lser 2 4 4.51086218E-10
C1 3 4 0.000000015
Rpar 3 4 6700000000
.ends 0805_885012207123_15nF
*******
.subckt 0805_885012207124_22nF 1 2
Rser 1 3 0.05
Lser 2 4 5.34340678E-10
C1 3 4 0.000000022
Rpar 3 4 4500000000
.ends 0805_885012207124_22nF
*******
.subckt 0805_885012207125_33nF 1 2
Rser 1 3 0.027855481442
Lser 2 4 4.0266816E-10
C1 3 4 0.000000033
Rpar 3 4 3000000000
.ends 0805_885012207125_33nF
*******
.subckt 0805_885012207126_47nF 1 2
Rser 1 3 0.0193681345947
Lser 2 4 3.56511593E-10
C1 3 4 0.000000047
Rpar 3 4 2100000000
.ends 0805_885012207126_47nF
*******
.subckt 0805_885012207127_68nF 1 2
Rser 1 3 0.0131992658565
Lser 2 4 3.66797021E-10
C1 3 4 0.000000068
Rpar 3 4 1500000000
.ends 0805_885012207127_68nF
*******
.subckt 0805_885012207128_100nF 1 2
Rser 1 3 0.0114794409661
Lser 2 4 3.71233852E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0805_885012207128_100nF
*******
.subckt 1206_885012208101_150pF 1 2
Rser 1 3 0.70365102611
Lser 2 4 3.78992769E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012208101_150pF
*******
.subckt 1206_885012208103_330pF 1 2
Rser 1 3 0.416289638796
Lser 2 4 4.89828253E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012208103_330pF
*******
.subckt 1206_885012208104_470pF 1 2
Rser 1 3 0.362109688542
Lser 2 4 4.01551911E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208104_470pF
*******
.subckt 1206_885012208105_680pF 1 2
Rser 1 3 0.332767276854
Lser 2 4 5.5598151E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012208105_680pF
*******
.subckt 1206_885012208106_1nF 1 2
Rser 1 3 0.24361864545
Lser 2 4 4.48764151E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208106_1nF
*******
.subckt 1206_885012208107_1.5nF 1 2
Rser 1 3 0.185507432166
Lser 2 4 4.5702585E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012208107_1.5nF
*******
.subckt 1206_885012208109_3.3nF 1 2
Rser 1 3 0.123971561911
Lser 2 4 4.87780525E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012208109_3.3nF
*******
.subckt 1206_885012208110_4.7nF 1 2
Rser 1 3 0.1
Lser 2 4 0.00000000049
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208110_4.7nF
*******
.subckt 1206_885012208111_6.8nF 1 2
Rser 1 3 0.0785959830702
Lser 2 4 5.43016322E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012208111_6.8nF
*******
.subckt 1206_885012208112_10nF 1 2
Rser 1 3 0.0821267479008
Lser 2 4 5.05894889E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208112_10nF
*******
.subckt 1206_885012208113_15nF 1 2
Rser 1 3 0.0562607370369
Lser 2 4 5.19798206E-10
C1 3 4 0.000000015
Rpar 3 4 6700000000
.ends 1206_885012208113_15nF
*******
.subckt 1206_885012208115_33nF 1 2
Rser 1 3 0.0633889215043
Lser 2 4 5.17142938E-10
C1 3 4 0.000000033
Rpar 3 4 3000000000
.ends 1206_885012208115_33nF
*******
.subckt 1206_885012208116_47nF 1 2
Rser 1 3 0.0362676531527
Lser 2 4 5.26289035E-10
C1 3 4 0.000000047
Rpar 3 4 2100000000
.ends 1206_885012208116_47nF
*******
.subckt 1206_885012208117_68nF 1 2
Rser 1 3 0.0206252921491
Lser 2 4 4.8689903E-10
C1 3 4 0.000000068
Rpar 3 4 1500000000
.ends 1206_885012208117_68nF
*******
.subckt 1206_885012208118_100nF 1 2
Rser 1 3 0.0147498855833
Lser 2 4 5.50636098E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1206_885012208118_100nF
*******
.subckt 1206_885012208119_150nF 1 2
Rser 1 3 0.00800974723287
Lser 2 4 3.65669763E-10
C1 3 4 0.00000015
Rpar 3 4 700000000
.ends 1206_885012208119_150nF
*******
.subckt 1210_885012209069_1uF 1 2
Rser 1 3 0.0053441098735
Lser 2 4 6.51295361E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 1210_885012209069_1uF
*******
.subckt 1210_885012209071_2.2uF 1 2
Rser 1 3 0.014
Lser 2 4 0.000000000755
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 1210_885012209071_2.2uF
*******
.subckt 2220_885012214001_10uF 1 2
Rser 1 3 0.003
Lser 2 4 0.0000000012
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 2220_885012214001_10uF
*******
.subckt 2220_885012214002_3.3uF 1 2
Rser 1 3 0.0056
Lser 2 4 0.0000000012
C1 3 4 0.0000033
Rpar 3 4 30000000
.ends 2220_885012214002_3.3uF
*******
.subckt 2220_885012214003_4.7uF 1 2
Rser 1 3 0.0043
Lser 2 4 0.0000000013
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 2220_885012214003_4.7uF
*******
.subckt 2220_885012214006_10uF 1 2
Rser 1 3 0.003
Lser 2 4 0.0000000012
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 2220_885012214006_10uF
*******
.subckt 0805_885012207130_470nF 1 2
Rser 1 3 0.011
Lser 2 4 0.0000000009
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0805_885012207130_470nF
*******
.subckt 0402_885012005020_1.5pF 1 2
Rser 1 3 1.045
Lser 2 4 0.00000000035
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0402_885012005020_1.5pF
*******
.subckt 0402_885012005021_2.2pF 1 2
Rser 1 3 0.37427104318
Lser 2 4 2.39727122E-10
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0402_885012005021_2.2pF
*******
.subckt 0402_885012005022_3.3pF 1 2
Rser 1 3 0.394048440694
Lser 2 4 2.60787564E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0402_885012005022_3.3pF
*******
.subckt 0402_885012005023_4.7pF 1 2
Rser 1 3 0.475944818481
Lser 2 4 2.97209578E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0402_885012005023_4.7pF
*******
.subckt 0402_885012005024_6.8pF 1 2
Rser 1 3 0.357812051681
Lser 2 4 2.43515953E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0402_885012005024_6.8pF
*******
.subckt 0402_885012005025_10pF 1 2
Rser 1 3 0.486385754904
Lser 2 4 3.42455186E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005025_10pF
*******
.subckt 0402_885012005026_15pF 1 2
Rser 1 3 0.385031326079
Lser 2 4 3.02592165E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885012005026_15pF
*******
.subckt 0402_885012005027_22pF 1 2
Rser 1 3 0.304814718575
Lser 2 4 3.0242914E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885012005027_22pF
*******
.subckt 0402_885012005028_33pF 1 2
Rser 1 3 0.244839252069
Lser 2 4 2.43449082E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005028_33pF
*******
.subckt 0402_885012005029_47pF 1 2
Rser 1 3 0.199232330322
Lser 2 4 2.79396057E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005029_47pF
*******
.subckt 0402_885012005030_68pF 1 2
Rser 1 3 0.183246570883
Lser 2 4 2.43281747E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005030_68pF
*******
.subckt 0402_885012005031_100pF 1 2
Rser 1 3 0.125698815083
Lser 2 4 2.36883012E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005031_100pF
*******
.subckt 0402_885012005032_150pF 1 2
Rser 1 3 0.0914737764723
Lser 2 4 2.04884984E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012005032_150pF
*******
.subckt 0402_885012005033_220pF 1 2
Rser 1 3 0.0784599744138
Lser 2 4 2.05801081E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012005033_220pF
*******
.subckt 0603_885012006017_10pF 1 2
Rser 1 3 0.4238423835
Lser 2 4 6.15454653E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006017_10pF
*******
.subckt 0603_885012006018_15pF 1 2
Rser 1 3 0.331903216145
Lser 2 4 4.69540847E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006018_15pF
*******
.subckt 0603_885012006019_22pF 1 2
Rser 1 3 0.348201721723
Lser 2 4 5.50963961E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006019_22pF
*******
.subckt 0603_885012006020_33pF 1 2
Rser 1 3 0.337785757957
Lser 2 4 7.34244223E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006020_33pF
*******
.subckt 0603_885012006021_47pF 1 2
Rser 1 3 0.256261040981
Lser 2 4 6.94150338E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006021_47pF
*******
.subckt 0603_885012006022_68pF 1 2
Rser 1 3 0.161913740901
Lser 2 4 6.38999674E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006022_68pF
*******
.subckt 0603_885012006023_100pF 1 2
Rser 1 3 0.123459009657
Lser 2 4 6.00573816E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006023_100pF
*******
.subckt 0603_885012006024_150pF 1 2
Rser 1 3 0.110788543459
Lser 2 4 5.59777275E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006024_150pF
*******
.subckt 0603_885012006025_220pF 1 2
Rser 1 3 0.0988385216426
Lser 2 4 5.64504761E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012006025_220pF
*******
.subckt 0603_885012006026_330pF 1 2
Rser 1 3 0.0877208643899
Lser 2 4 5.53240043E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006026_330pF
*******
.subckt 0603_885012006027_470pF 1 2
Rser 1 3 0.0602974058901
Lser 2 4 5.48330767E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006027_470pF
*******
.subckt 0603_885012006028_680pF 1 2
Rser 1 3 0.0523826835624
Lser 2 4 5.05789539E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006028_680pF
*******
.subckt 0603_885012006029_1nF 1 2
Rser 1 3 0.0440182000352
Lser 2 4 4.19702079E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006029_1nF
*******
.subckt 0805_885012007010_10pF 1 2
Rser 1 3 0.372486331807
Lser 2 4 3.46703717E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0805_885012007010_10pF
*******
.subckt 0805_885012007011_15pF 1 2
Rser 1 3 0.299277635225
Lser 2 4 4.59074821E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007011_15pF
*******
.subckt 0805_885012007012_22pF 1 2
Rser 1 3 0.353164620745
Lser 2 4 4.83956508E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0805_885012007012_22pF
*******
.subckt 0805_885012007013_33pF 1 2
Rser 1 3 0.253567178585
Lser 2 4 4.67181086E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007013_33pF
*******
.subckt 0805_885012007014_47pF 1 2
Rser 1 3 0.224186907869
Lser 2 4 4.55318299E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885012007014_47pF
*******
.subckt 0805_885012007015_68pF 1 2
Rser 1 3 0.177556084991
Lser 2 4 3.40488342E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0805_885012007015_68pF
*******
.subckt 0805_885012007016_100pF 1 2
Rser 1 3 0.144693224126
Lser 2 4 2.25885151E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007016_100pF
*******
.subckt 0805_885012007017_150pF 1 2
Rser 1 3 0.123365902974
Lser 2 4 2.19751744E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007017_150pF
*******
.subckt 0805_885012007018_220pF 1 2
Rser 1 3 0.10837087132
Lser 2 4 2.252525E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012007018_220pF
*******
.subckt 0805_885012007019_330pF 1 2
Rser 1 3 0.0921576071204
Lser 2 4 2.40260993E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007019_330pF
*******
.subckt 0805_885012007020_470pF 1 2
Rser 1 3 0.0750834191209
Lser 2 4 2.93018556E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007020_470pF
*******
.subckt 0805_885012007021_1nF 1 2
Rser 1 3 0.0483999213452
Lser 2 4 2.79211981E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007021_1nF
*******
.subckt 0805_885012007022_1.5nF 1 2
Rser 1 3 0.0373928905809
Lser 2 4 2.95075489E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012007022_1.5nF
*******
.subckt 0805_885012007023_2.2nF 1 2
Rser 1 3 0.0368859488683
Lser 2 4 2.79156194E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012007023_2.2nF
*******
.subckt 0805_885012007024_3.3nF 1 2
Rser 1 3 0.0117602115678
Lser 2 4 2.50664287E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012007024_3.3nF
*******
.subckt 0805_885012007025_4.7nF 1 2
Rser 1 3 0.0198836793746
Lser 2 4 1.51240813E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012007025_4.7nF
*******
.subckt 1206_885012008011_22pF 1 2
Rser 1 3 0.324375840883
Lser 2 4 5.44232375E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1206_885012008011_22pF
*******
.subckt 1206_885012008012_100pF 1 2
Rser 1 3 0.141237836467
Lser 2 4 5.16904289E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008012_100pF
*******
.subckt 1206_885012008013_150pF 1 2
Rser 1 3 0.123922377922
Lser 2 4 4.91328479E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012008013_150pF
*******
.subckt 1206_885012008014_220pF 1 2
Rser 1 3 0.0914487723967
Lser 2 4 4.26746797E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012008014_220pF
*******
.subckt 1206_885012008015_2.2nF 1 2
Rser 1 3 0.0540944991554
Lser 2 4 4.14167967E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012008015_2.2nF
*******
.subckt 1206_885012008016_6.8nF 1 2
Rser 1 3 0.0272311989762
Lser 2 4 3.46260293E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008016_6.8nF
*******
.subckt 1206_885012008017_10nF 1 2
Rser 1 3 0.0157731913832
Lser 2 4 3.49723643E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008017_10nF
*******
.subckt 1210_885012009001_15nF 1 2
Rser 1 3 0.0355230024751
Lser 2 4 8.2968558E-11
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1210_885012009001_15nF
*******
.subckt 1812_885012010001_1nF 1 2
Rser 1 3 0.0510603999373
Lser 2 4 2.97374009E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_885012010001_1nF
*******
.subckt 1812_885012010002_22nF 1 2
Rser 1 3 0.0138901707005
Lser 2 4 3.25297738E-10
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1812_885012010002_22nF
*******
.subckt 0402_885012105014_33nF 1 2
Rser 1 3 0.026490919016
Lser 2 4 2.00303378E-10
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0402_885012105014_33nF
*******
.subckt 0402_885012105015_47nF 1 2
Rser 1 3 0.0367849496471
Lser 2 4 1.808767E-10
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0402_885012105015_47nF
*******
.subckt 0402_885012105016_100nF 1 2
Rser 1 3 0.018877276336
Lser 2 4 3.14688963E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012105016_100nF
*******
.subckt 0402_885012105017_220nF 1 2
Rser 1 3 0.0118013539585
Lser 2 4 3.47460059E-10
C1 3 4 0.00000022
Rpar 3 4 500000000
.ends 0402_885012105017_220nF
*******
.subckt 0603_885012106013_220nF 1 2
Rser 1 3 0.0111678211386
Lser 2 4 2.40956055E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012106013_220nF
*******
.subckt 0603_885012106014_330nF 1 2
Rser 1 3 0.0117435280097
Lser 2 4 3.10748007E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012106014_330nF
*******
.subckt 0603_885012106015_470nF 1 2
Rser 1 3 0.0117435280097
Lser 2 4 2.50748007E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012106015_470nF
*******
.subckt 0603_885012106016_680nF 1 2
Rser 1 3 0.0127619086118
Lser 2 4 3.65801201E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0603_885012106016_680nF
*******
.subckt 0603_885012106017_1uF 1 2
Rser 1 3 0.00745135412008
Lser 2 4 3.04086627E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012106017_1uF
*******
.subckt 0603_885012106018_2.2uF 1 2
Rser 1 3 0.00721183501635
Lser 2 4 2.59345303E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0603_885012106018_2.2uF
*******
.subckt 0805_885012107012_2.2uF 1 2
Rser 1 3 0.0046352610288
Lser 2 4 2.55261723E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012107012_2.2uF
*******
.subckt 0805_885012107013_4.7uF 1 2
Rser 1 3 0.0035599941357
Lser 2 4 2.56410699E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0805_885012107013_4.7uF
*******
.subckt 0805_885012107014_10uF 1 2
Rser 1 3 0.0034022396539
Lser 2 4 3.00259834E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0805_885012107014_10uF
*******
.subckt 1206_885012108013_1.5uF 1 2
Rser 1 3 0.0096965404251
Lser 2 4 6.58515557E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 1206_885012108013_1.5uF
*******
.subckt 1206_885012108014_2.2uF 1 2
Rser 1 3 0.00698767716064
Lser 2 4 5.83531315E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012108014_2.2uF
*******
.subckt 1206_885012108015_3.3uF 1 2
Rser 1 3 0.00545085791999
Lser 2 4 6.21772385E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012108015_3.3uF
*******
.subckt 1206_885012108016_4.7uF 1 2
Rser 1 3 0.00700055770575
Lser 2 4 5.37514029E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1206_885012108016_4.7uF
*******
.subckt 1206_885012108017_10uF 1 2
Rser 1 3 0.00377815297038
Lser 2 4 8.77331047E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1206_885012108017_10uF
*******
.subckt 1206_885012108018_22uF 1 2
Rser 1 3 0.00326232270901
Lser 2 4 5.38545474E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1206_885012108018_22uF
*******
.subckt 1210_885012109008_4.7uF 1 2
Rser 1 3 0.0035836083267
Lser 2 4 3.35721238E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012109008_4.7uF
*******
.subckt 1210_885012109009_10uF 1 2
Rser 1 3 0.00244609668461
Lser 2 4 7.73879687E-10
C1 3 4 0.00001
Rpar 3 4 50000000
.ends 1210_885012109009_10uF
*******
.subckt 1210_885012109010_22uF 1 2
Rser 1 3 0.00405759674222
Lser 2 4 1.477484223E-09
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1210_885012109010_22uF
*******
.subckt 1210_885012109011_47uF 1 2
Rser 1 3 0.00225907860771
Lser 2 4 0.0000000009
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1210_885012109011_47uF
*******
.subckt 0402_885012205019_100pF 1 2
Rser 1 3 0.77428
Lser 2 4 0.00000000014154
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012205019_100pF
*******
.subckt 0402_885012205020_150pF 1 2
Rser 1 3 0.67192
Lser 2 4 0.00000000015134
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012205020_150pF
*******
.subckt 0402_885012205021_220pF 1 2
Rser 1 3 0.5734
Lser 2 4 0.00000000018579
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012205021_220pF
*******
.subckt 0402_885012205022_330pF 1 2
Rser 1 3 0.41636
Lser 2 4 0.000000000183
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012205022_330pF
*******
.subckt 0402_885012205023_470pF 1 2
Rser 1 3 0.31598
Lser 2 4 0.0000000002154
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012205023_470pF
*******
.subckt 0402_885012205024_680pF 1 2
Rser 1 3 0.23994
Lser 2 4 0.00000000014784
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0402_885012205024_680pF
*******
.subckt 0402_885012205025_1nF 1 2
Rser 1 3 0.213522308242
Lser 2 4 2.15925639E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205025_1nF
*******
.subckt 0402_885012205026_1.5nF 1 2
Rser 1 3 0.17301
Lser 2 4 0.00000000025499
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0402_885012205026_1.5nF
*******
.subckt 0402_885012205027_2.2nF 1 2
Rser 1 3 0.12141
Lser 2 4 0.00000000025109
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0402_885012205027_2.2nF
*******
.subckt 0402_885012205028_3.3nF 1 2
Rser 1 3 0.08715
Lser 2 4 0.00000000022723
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0402_885012205028_3.3nF
*******
.subckt 0402_885012205029_4.7nF 1 2
Rser 1 3 0.07998
Lser 2 4 0.00000000017442
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205029_4.7nF
*******
.subckt 0402_885012205030_6.8nF 1 2
Rser 1 3 0.07283
Lser 2 4 0.00000000019034
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0402_885012205030_6.8nF
*******
.subckt 0402_885012205031_10nF 1 2
Rser 1 3 0.05542
Lser 2 4 0.00000000019893
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0402_885012205031_10nF
*******
.subckt 0402_885012205032_15nF 1 2
Rser 1 3 0.04045
Lser 2 4 0.00000000020744
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0402_885012205032_15nF
*******
.subckt 0402_885012205033_22nF 1 2
Rser 1 3 0.02779
Lser 2 4 0.00000000018757
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0402_885012205033_22nF
*******
.subckt 0402_885012205034_33nF 1 2
Rser 1 3 0.01627
Lser 2 4 0.00000000021013
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0402_885012205034_33nF
*******
.subckt 0402_885012205035_47nF 1 2
Rser 1 3 0.0085
Lser 2 4 0.00000000020707
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0402_885012205035_47nF
*******
.subckt 0402_885012205036_68nF 1 2
Rser 1 3 0.01842
Lser 2 4 0.00000000022333
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0402_885012205036_68nF
*******
.subckt 0402_885012205037_100nF 1 2
Rser 1 3 0.0169137492565
Lser 2 4 3.31963015E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205037_100nF
*******
.subckt 0402_885012205037R_100nF 1 2
Rser 1 3 0.0169137492565
Lser 2 4 3.31963015E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205037R_100nF
*******
.subckt 0603_885012206028_100pF 1 2
Rser 1 3 0.83279
Lser 2 4 0.00000000026283
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206028_100pF
*******
.subckt 0603_885012206029_150pF 1 2
Rser 1 3 0.68443
Lser 2 4 0.00000000029041
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012206029_150pF
*******
.subckt 0603_885012206030_220pF 1 2
Rser 1 3 0.49382
Lser 2 4 0.00000000028774
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012206030_220pF
*******
.subckt 0603_885012206031_330pF 1 2
Rser 1 3 0.4404
Lser 2 4 0.00000000034035
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206031_330pF
*******
.subckt 0603_885012206032_470pF 1 2
Rser 1 3 0.32027
Lser 2 4 0.00000000032279
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206032_470pF
*******
.subckt 0603_885012206033_680pF 1 2
Rser 1 3 0.31076
Lser 2 4 0.00000000037089
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206033_680pF
*******
.subckt 0603_885012206034_1nF 1 2
Rser 1 3 0.2266
Lser 2 4 0.00000000040041
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206034_1nF
*******
.subckt 0603_885012206035_1.5nF 1 2
Rser 1 3 0.13944
Lser 2 4 0.00000000032692
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206035_1.5nF
*******
.subckt 0603_885012206036_2.2nF 1 2
Rser 1 3 0.12185
Lser 2 4 0.00000000030888
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012206036_2.2nF
*******
.subckt 0603_885012206037_3.3nF 1 2
Rser 1 3 0.0993
Lser 2 4 0.00000000030024
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206037_3.3nF
*******
.subckt 0603_885012206038_4.7nF 1 2
Rser 1 3 0.0825557398709
Lser 2 4 2.58966471E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206038_4.7nF
*******
.subckt 0603_885012206039_6.8nF 1 2
Rser 1 3 0.06147
Lser 2 4 0.00000000035083
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206039_6.8nF
*******
.subckt 0603_885012206040_10nF 1 2
Rser 1 3 0.06145
Lser 2 4 0.00000000036058
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206040_10nF
*******
.subckt 0603_885012206041_15nF 1 2
Rser 1 3 0.04438
Lser 2 4 0.00000000031844
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0603_885012206041_15nF
*******
.subckt 0603_885012206042_22nF 1 2
Rser 1 3 0.03181
Lser 2 4 0.00000000024225
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885012206042_22nF
*******
.subckt 0603_885012206043_33nF 1 2
Rser 1 3 0.02195
Lser 2 4 0.00000000030558
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0603_885012206043_33nF
*******
.subckt 0603_885012206044_47nF 1 2
Rser 1 3 0.01525
Lser 2 4 0.00000000027141
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0603_885012206044_47nF
*******
.subckt 0603_885012206045_68nF 1 2
Rser 1 3 0.01508
Lser 2 4 0.00000000030779
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0603_885012206045_68nF
*******
.subckt 0603_885012206046_100nF 1 2
Rser 1 3 0.0189313024822
Lser 2 4 4.50736859E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206046_100nF
*******
.subckt 0603_885012206047_150nF 1 2
Rser 1 3 0.0192205094865
Lser 2 4 4.7670705E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0603_885012206047_150nF
*******
.subckt 0603_885012206048_220nF 1 2
Rser 1 3 0.0139027111992
Lser 2 4 4.40984618E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012206048_220nF
*******
.subckt 0603_885012206049_330nF 1 2
Rser 1 3 0.0117878976558
Lser 2 4 3.9313295E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012206049_330nF
*******
.subckt 0603_885012206050_470nF 1 2
Rser 1 3 0.00930503966198
Lser 2 4 4.27988831E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012206050_470nF
*******
.subckt 0603_885012206051_680nF 1 2
Rser 1 3 0.00730097281816
Lser 2 4 4.2920775E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0603_885012206051_680nF
*******
.subckt 0603_885012206052_1uF 1 2
Rser 1 3 0.00742821402486
Lser 2 4 2.51142993E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012206052_1uF
*******
.subckt 0805_885012207027_100pF 1 2
Rser 1 3 0.8158
Lser 2 4 0.00000000024681
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207027_100pF
*******
.subckt 0805_885012207028_150pF 1 2
Rser 1 3 0.69537
Lser 2 4 0.00000000030323
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012207028_150pF
*******
.subckt 0805_885012207029_220pF 1 2
Rser 1 3 0.49653
Lser 2 4 0.00000000027715
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012207029_220pF
*******
.subckt 0805_885012207030_330pF 1 2
Rser 1 3 0.28432
Lser 2 4 0.00000000020282
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012207030_330pF
*******
.subckt 0805_885012207031_470pF 1 2
Rser 1 3 0.19262
Lser 2 4 0.00000000022289
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207031_470pF
*******
.subckt 0805_885012207032_680pF 1 2
Rser 1 3 0.15908
Lser 2 4 0.00000000028074
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012207032_680pF
*******
.subckt 0805_885012207033_1nF 1 2
Rser 1 3 0.10327
Lser 2 4 0.00000000021794
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207033_1nF
*******
.subckt 0805_885012207034_1.5nF 1 2
Rser 1 3 0.0607
Lser 2 4 0.00000000029167
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207034_1.5nF
*******
.subckt 0805_885012207035_2.2nF 1 2
Rser 1 3 0.0294
Lser 2 4 0.00000000027896
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012207035_2.2nF
*******
.subckt 0805_885012207036_3.3nF 1 2
Rser 1 3 0.00336
Lser 2 4 0.00000000024965
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207036_3.3nF
*******
.subckt 0805_885012207037_4.7nF 1 2
Rser 1 3 0.02846
Lser 2 4 0.00000000015236
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012207037_4.7nF
*******
.subckt 0805_885012207038_6.8nF 1 2
Rser 1 3 0.07854
Lser 2 4 0.00000000032137
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0805_885012207038_6.8nF
*******
.subckt 0805_885012207039_10nF 1 2
Rser 1 3 0.06279
Lser 2 4 0.00000000033683
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207039_10nF
*******
.subckt 0805_885012207040_15nF 1 2
Rser 1 3 0.05886
Lser 2 4 0.000000000349367
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0805_885012207040_15nF
*******
.subckt 0805_885012207041_22nF 1 2
Rser 1 3 0.04639
Lser 2 4 0.00000000031523
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0805_885012207041_22nF
*******
.subckt 0805_885012207042_33nF 1 2
Rser 1 3 0.03915
Lser 2 4 0.0000000003028
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0805_885012207042_33nF
*******
.subckt 0805_885012207043_47nF 1 2
Rser 1 3 0.04259
Lser 2 4 0.000000000307
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0805_885012207043_47nF
*******
.subckt 0805_885012207044_68nF 1 2
Rser 1 3 0.02591
Lser 2 4 0.00000000028743
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0805_885012207044_68nF
*******
.subckt 0805_885012207045_100nF 1 2
Rser 1 3 0.0170178433002
Lser 2 4 0.00000000038
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207045_100nF
*******
.subckt 0805_885012207046_150nF 1 2
Rser 1 3 0.0131969599932
Lser 2 4 4.43917137E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0805_885012207046_150nF
*******
.subckt 0805_885012207047_220nF 1 2
Rser 1 3 0.0124886466337
Lser 2 4 0.0000000003
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885012207047_220nF
*******
.subckt 0805_885012207048_330nF 1 2
Rser 1 3 0.0121631731335
Lser 2 4 0.00000000036
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885012207048_330nF
*******
.subckt 0805_885012207049_470nF 1 2
Rser 1 3 0.00820167627427
Lser 2 4 0.00000000049
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0805_885012207049_470nF
*******
.subckt 0805_885012207050_680nF 1 2
Rser 1 3 0.00778029663502
Lser 2 4 0.000000000512
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0805_885012207050_680nF
*******
.subckt 0805_885012207051_1uF 1 2
Rser 1 3 0.0071335712548
Lser 2 4 2.56885128E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885012207051_1uF
*******
.subckt 0805_885012207052_2.2uF 1 2
Rser 1 3 0.00474724521779
Lser 2 4 2.59969084E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012207052_2.2uF
*******
.subckt 0805_885012207053_4.7uF 1 2
Rser 1 3 0.00357806469138
Lser 2 4 4.01525773E-10
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0805_885012207053_4.7uF
*******
.subckt 1206_885012208020_220pF 1 2
Rser 1 3 0.54413
Lser 2 4 0.00000000031019
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012208020_220pF
*******
.subckt 1206_885012208021_470pF 1 2
Rser 1 3 0.34
Lser 2 4 0.00000000042098
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208021_470pF
*******
.subckt 1206_885012208022_1nF 1 2
Rser 1 3 0.23809
Lser 2 4 0.00000000043011
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208022_1nF
*******
.subckt 1206_885012208023_2.2nF 1 2
Rser 1 3 0.16161
Lser 2 4 0.0000000004207
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012208023_2.2nF
*******
.subckt 1206_885012208024_3.3nF 1 2
Rser 1 3 0.12067
Lser 2 4 0.00000000046077
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012208024_3.3nF
*******
.subckt 1206_885012208025_4.7nF 1 2
Rser 1 3 0.1467
Lser 2 4 0.00000000046584
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208025_4.7nF
*******
.subckt 1206_885012208026_10nF 1 2
Rser 1 3 0.07047
Lser 2 4 0.0000000006906
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208026_10nF
*******
.subckt 1206_885012208027_22nF 1 2
Rser 1 3 0.05191
Lser 2 4 0.00000000044884
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1206_885012208027_22nF
*******
.subckt 1206_885012208028_33nF 1 2
Rser 1 3 0.05461
Lser 2 4 0.00000000071542
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1206_885012208028_33nF
*******
.subckt 1206_885012208029_47nF 1 2
Rser 1 3 0.0511
Lser 2 4 0.00000000044681
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1206_885012208029_47nF
*******
.subckt 1206_885012208030_100nF 1 2
Rser 1 3 0.0236394219015
Lser 2 4 6.65660931E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885012208030_100nF
*******
.subckt 1206_885012208031_150nF 1 2
Rser 1 3 0.0172296802581
Lser 2 4 6.75934228E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1206_885012208031_150nF
*******
.subckt 1206_885012208032_220nF 1 2
Rser 1 3 0.0123092011142
Lser 2 4 6.56591189E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1206_885012208032_220nF
*******
.subckt 1206_885012208033_330nF 1 2
Rser 1 3 0.0121092486479
Lser 2 4 7.02655219E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1206_885012208033_330nF
*******
.subckt 1206_885012208034_470nF 1 2
Rser 1 3 0.0106020491014
Lser 2 4 7.42809674E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1206_885012208034_470nF
*******
.subckt 1206_885012208035_680nF 1 2
Rser 1 3 0.00686375950243
Lser 2 4 7.21249479E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1206_885012208035_680nF
*******
.subckt 1206_885012208036_1uF 1 2
Rser 1 3 0.00696547352182
Lser 2 4 6.33927755E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885012208036_1uF
*******
.subckt 1206_885012208037_1.5uF 1 2
Rser 1 3 0.00838199168584
Lser 2 4 6.76254119E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 1206_885012208037_1.5uF
*******
.subckt 1206_885012208038_2.2uF 1 2
Rser 1 3 0.00657322849514
Lser 2 4 5.35127467E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012208038_2.2uF
*******
.subckt 1206_885012208039_3.3uF 1 2
Rser 1 3 0.00583502254442
Lser 2 4 5.58875803E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012208039_3.3uF
*******
.subckt 1206_885012208040_4.7uF 1 2
Rser 1 3 0.00382284206604
Lser 2 4 7.81956777E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1206_885012208040_4.7uF
*******
.subckt 1206_885012208041_10uF 1 2
Rser 1 3 0.00303
Lser 2 4 0.00000000078818
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1206_885012208041_10uF
*******
.subckt 1210_885012209007_150nF 1 2
Rser 1 3 0.0143454209584
Lser 2 4 5.36188212E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1210_885012209007_150nF
*******
.subckt 1210_885012209008_220nF 1 2
Rser 1 3 0.01034976783
Lser 2 4 5.13522247E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1210_885012209008_220nF
*******
.subckt 1210_885012209009_470nF 1 2
Rser 1 3 0.00837032621271
Lser 2 4 5.45617858E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1210_885012209009_470nF
*******
.subckt 1210_885012209010_680nF 1 2
Rser 1 3 0.00546743874253
Lser 2 4 5.62694253E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1210_885012209010_680nF
*******
.subckt 1210_885012209011_1uF 1 2
Rser 1 3 0.00410122631789
Lser 2 4 3.71398434E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209011_1uF
*******
.subckt 1210_885012209012_2.2uF 1 2
Rser 1 3 0.0039891272832
Lser 2 4 5.25018615E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1210_885012209012_2.2uF
*******
.subckt 1210_885012209013_4.7uF 1 2
Rser 1 3 0.00524566546715
Lser 2 4 5.20085349E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012209013_4.7uF
*******
.subckt 1210_885012209014_10uF 1 2
Rser 1 3 0.00222604043193
Lser 2 4 7.58236705E-10
C1 3 4 0.00001
Rpar 3 4 100000000
.ends 1210_885012209014_10uF
*******
.subckt 1812_885012210001_10nF 1 2
Rser 1 3 0.07465
Lser 2 4 0.00000000052475
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012210001_10nF
*******
.subckt 1812_885012210002_47nF 1 2
Rser 1 3 0.03429
Lser 2 4 0.00000000074448
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1812_885012210002_47nF
*******
.subckt 1812_885012210003_680nF 1 2
Rser 1 3 0.00789799680346
Lser 2 4 5.51300911E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1812_885012210003_680nF
*******
.subckt 1812_885012210004_1uF 1 2
Rser 1 3 0.00726915726357
Lser 2 4 3.95869894E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1812_885012210004_1uF
*******
.subckt 0201_885012104001_100nF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000008
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0201_885012104001_100nF
*******
.subckt 0201_885012104007_1uF 1 2
Rser 1 3 0.01366
Lser 2 4 0.000000000165
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0201_885012104007_1uF
*******
.subckt 0603_885012106029_2.2uF 1 2
Rser 1 3 0.011
Lser 2 4 0.0000000008
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0603_885012106029_2.2uF
*******
.subckt 0402_885012005034_1pF 1 2
Rser 1 3 0.734
Lser 2 4 0.00000000038
C1 3 4 0.000000000001
Rpar 3 4 10000000000
.ends 0402_885012005034_1pF
*******
.subckt 0402_885012005040_10pF 1 2
Rser 1 3 0.467848447943
Lser 2 4 3.77046381E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005040_10pF
*******
.subckt 0402_885012005041_15pF 1 2
Rser 1 3 0.34552139712
Lser 2 4 3.31461104E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885012005041_15pF
*******
.subckt 0402_885012005042_22pF 1 2
Rser 1 3 0.285282706764
Lser 2 4 3.08207076E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885012005042_22pF
*******
.subckt 0402_885012005043_33pF 1 2
Rser 1 3 0.230231956882
Lser 2 4 2.96875149E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005043_33pF
*******
.subckt 0402_885012005044_47pF 1 2
Rser 1 3 0.203455175683
Lser 2 4 3.46537476E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005044_47pF
*******
.subckt 0402_885012005045_68pF 1 2
Rser 1 3 0.18781473697
Lser 2 4 3.22027908E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005045_68pF
*******
.subckt 0402_885012005046_100pF 1 2
Rser 1 3 0.0759217345208
Lser 2 4 3.94922966E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005046_100pF
*******
.subckt 0402_885012005047_150pF 1 2
Rser 1 3 0.112246046138
Lser 2 4 2.15549473E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012005047_150pF
*******
.subckt 0402_885012005048_220pF 1 2
Rser 1 3 0.104232515193
Lser 2 4 1.92172989E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012005048_220pF
*******
.subckt 0603_885012006030_4.7pF 1 2
Rser 1 3 0.29124727578
Lser 2 4 4.29705418E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0603_885012006030_4.7pF
*******
.subckt 0603_885012006031_6.8pF 1 2
Rser 1 3 0.299024437013
Lser 2 4 4.5809474E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0603_885012006031_6.8pF
*******
.subckt 0603_885012006032_10pF 1 2
Rser 1 3 0.445774201336
Lser 2 4 4.28073844E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006032_10pF
*******
.subckt 0603_885012006033_15pF 1 2
Rser 1 3 0.353119905486
Lser 2 4 4.35266975E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006033_15pF
*******
.subckt 0603_885012006034_22pF 1 2
Rser 1 3 0.352481322316
Lser 2 4 5.8820344E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006034_22pF
*******
.subckt 0603_885012006035_33pF 1 2
Rser 1 3 0.305919966941
Lser 2 4 5.25713034E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006035_33pF
*******
.subckt 0603_885012006036_47pF 1 2
Rser 1 3 0.062255914612
Lser 2 4 4.24328623E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006036_47pF
*******
.subckt 0603_885012006037_68pF 1 2
Rser 1 3 0.159672910297
Lser 2 4 6.46220787E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006037_68pF
*******
.subckt 0603_885012006038_100pF 1 2
Rser 1 3 0.130130495234
Lser 2 4 5.8979323E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006038_100pF
*******
.subckt 0603_885012006039_150pF 1 2
Rser 1 3 0.097154893647
Lser 2 4 5.82598828E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006039_150pF
*******
.subckt 0603_885012006040_220pF 1 2
Rser 1 3 0.111748485631
Lser 2 4 6.02628009E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012006040_220pF
*******
.subckt 0603_885012006041_330pF 1 2
Rser 1 3 0.0829140919635
Lser 2 4 3.85173897E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006041_330pF
*******
.subckt 0603_885012006042_470pF 1 2
Rser 1 3 0.0647178553788
Lser 2 4 3.67931779E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006042_470pF
*******
.subckt 0603_885012006043_680pF 1 2
Rser 1 3 0.0641029132415
Lser 2 4 3.05763584E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006043_680pF
*******
.subckt 0603_885012006044_1nF 1 2
Rser 1 3 0.0419451701409
Lser 2 4 4.48170961E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006044_1nF
*******
.subckt 0805_885012007026_3.3pF 1 2
Rser 1 3 0.407676004204
Lser 2 4 4.49191488E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0805_885012007026_3.3pF
*******
.subckt 0805_885012007027_6.8pF 1 2
Rser 1 3 0.359480200218
Lser 2 4 4.5722648E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0805_885012007027_6.8pF
*******
.subckt 0805_885012007028_10pF 1 2
Rser 1 3 0.366485482781
Lser 2 4 5.23706793E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0805_885012007028_10pF
*******
.subckt 0805_885012007029_15pF 1 2
Rser 1 3 0.322140605571
Lser 2 4 5.33099942E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007029_15pF
*******
.subckt 0805_885012007030_22pF 1 2
Rser 1 3 0.337501541959
Lser 2 4 6.08362599E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0805_885012007030_22pF
*******
.subckt 0805_885012007031_33pF 1 2
Rser 1 3 0.266905660637
Lser 2 4 5.7081292E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007031_33pF
*******
.subckt 0805_885012007032_47pF 1 2
Rser 1 3 0.224971777912
Lser 2 4 5.50463607E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885012007032_47pF
*******
.subckt 0805_885012007033_68pF 1 2
Rser 1 3 0.188385732986
Lser 2 4 4.4496757E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0805_885012007033_68pF
*******
.subckt 0805_885012007034_100pF 1 2
Rser 1 3 0.118679326168
Lser 2 4 2.41991847E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007034_100pF
*******
.subckt 0805_885012007035_150pF 1 2
Rser 1 3 0.135556605699
Lser 2 4 4.3127146E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007035_150pF
*******
.subckt 0805_885012007036_220pF 1 2
Rser 1 3 0.115723179071
Lser 2 4 4.36175568E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012007036_220pF
*******
.subckt 0805_885012007037_330pF 1 2
Rser 1 3 0.0911424032195
Lser 2 4 4.34684674E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007037_330pF
*******
.subckt 0805_885012007038_470pF 1 2
Rser 1 3 0.0888157768288
Lser 2 4 4.59255914E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007038_470pF
*******
.subckt 0805_885012007039_680pF 1 2
Rser 1 3 0.0750121415022
Lser 2 4 4.46094349E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012007039_680pF
*******
.subckt 0805_885012007040_1nF 1 2
Rser 1 3 0.0506576337129
Lser 2 4 2.60606775E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007040_1nF
*******
.subckt 0805_885012007041_1.5nF 1 2
Rser 1 3 0.0403337213614
Lser 2 4 2.897145E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012007041_1.5nF
*******
.subckt 0805_885012007042_2.2nF 1 2
Rser 1 3 0.0313104040283
Lser 2 4 2.67647833E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012007042_2.2nF
*******
.subckt 0805_885012007043_3.3nF 1 2
Rser 1 3 0.0278586078187
Lser 2 4 3.06758727E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012007043_3.3nF
*******
.subckt 0805_885012007044_4.7nF 1 2
Rser 1 3 0.0125481242528
Lser 2 4 1.0825546E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012007044_4.7nF
*******
.subckt 1206_885012008019_10pF 1 2
Rser 1 3 0.391301643484
Lser 2 4 5.83813577E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1206_885012008019_10pF
*******
.subckt 1206_885012008020_33pF 1 2
Rser 1 3 0.254333105283
Lser 2 4 4.78321618E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 1206_885012008020_33pF
*******
.subckt 1206_885012008021_47pF 1 2
Rser 1 3 0.233708673806
Lser 2 4 4.88472845E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885012008021_47pF
*******
.subckt 1206_885012008022_68pF 1 2
Rser 1 3 0.199591933016
Lser 2 4 4.68378192E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 1206_885012008022_68pF
*******
.subckt 1206_885012008023_100pF 1 2
Rser 1 3 0.15525411437
Lser 2 4 4.47352225E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008023_100pF
*******
.subckt 1206_885012008024_330pF 1 2
Rser 1 3 0.0916318679708
Lser 2 4 3.11969377E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012008024_330pF
*******
.subckt 1206_885012008025_470pF 1 2
Rser 1 3 0.106551883888
Lser 2 4 4.30008474E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012008025_470pF
*******
.subckt 1206_885012008026_1nF 1 2
Rser 1 3 0.0693861515837
Lser 2 4 4.13253027E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012008026_1nF
*******
.subckt 1206_885012008027_2.2nF 1 2
Rser 1 3 0.0393800076857
Lser 2 4 5.03985839E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012008027_2.2nF
*******
.subckt 1206_885012008028_4.7nF 1 2
Rser 1 3 0.0260664466932
Lser 2 4 4.4983761E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012008028_4.7nF
*******
.subckt 1206_885012008029_6.8nF 1 2
Rser 1 3 0.0469294057584
Lser 2 4 4.43201944E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008029_6.8nF
*******
.subckt 1206_885012008030_10nF 1 2
Rser 1 3 0.0261734331747
Lser 2 4 5.33952576E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008030_10nF
*******
.subckt 1210_885012009002_1nF 1 2
Rser 1 3 0.0526199422099
Lser 2 4 2.28139939E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885012009002_1nF
*******
.subckt 1210_885012009003_2.2nF 1 2
Rser 1 3 0.236239384732
Lser 2 4 2.48857755E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1210_885012009003_2.2nF
*******
.subckt 1210_885012009004_4.7nF 1 2
Rser 1 3 0.0889145917519
Lser 2 4 2.66275966E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1210_885012009004_4.7nF
*******
.subckt 1210_885012009005_6.8nF 1 2
Rser 1 3 0.0165690812867
Lser 2 4 2.56210234E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1210_885012009005_6.8nF
*******
.subckt 1210_885012009006_15nF 1 2
Rser 1 3 0.0164446208365
Lser 2 4 3.024777E-10
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1210_885012009006_15nF
*******
.subckt 1812_885012010003_10nF 1 2
Rser 1 3 0.035610362113
Lser 2 4 2.40113972E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012010003_10nF
*******
.subckt 1812_885012010004_33nF 1 2
Rser 1 3 0.0120609525555
Lser 2 4 3.8469537E-10
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1812_885012010004_33nF
*******
.subckt 0402_885012105018_100nF 1 2
Rser 1 3 0.026120802334
Lser 2 4 3.09671131E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012105018_100nF
*******
.subckt 0603_885012106019_220nF 1 2
Rser 1 3 0.0108961182185
Lser 2 4 2.50789051E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012106019_220nF
*******
.subckt 0603_885012106020_470nF 1 2
Rser 1 3 0.00976845934589
Lser 2 4 2.50682976E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012106020_470nF
*******
.subckt 0603_885012106021_680nF 1 2
Rser 1 3 0.00991319698945
Lser 2 4 3.55175418E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0603_885012106021_680nF
*******
.subckt 0603_885012106022_1uF 1 2
Rser 1 3 0.00857861035867
Lser 2 4 3.03497279E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0603_885012106022_1uF
*******
.subckt 0603_885012106031_10uF 1 2
Rser 1 3 0.0105
Lser 2 4 0.0000000008
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 0603_885012106031_10uF
*******
.subckt 0805_885012107015_1uF 1 2
Rser 1 3 0.00799934804354
Lser 2 4 2.55135429E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885012107015_1uF
*******
.subckt 0805_885012107016_2.2uF 1 2
Rser 1 3 0.00497944150425
Lser 2 4 2.69972955E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012107016_2.2uF
*******
.subckt 0805_885012107017_3.3uF 1 2
Rser 1 3 0.0041415980008
Lser 2 4 2.72087954E-10
C1 3 4 0.0000033
Rpar 3 4 30000000
.ends 0805_885012107017_3.3uF
*******
.subckt 0805_885012107018_4.7uF 1 2
Rser 1 3 0.00349429730952
Lser 2 4 2.52123218E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0805_885012107018_4.7uF
*******
.subckt 1206_885012108019_2.2uF 1 2
Rser 1 3 0.00474329771021
Lser 2 4 5.16937352E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012108019_2.2uF
*******
.subckt 1206_885012108020_4.7uF 1 2
Rser 1 3 0.00541345635951
Lser 2 4 5.0768239E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1206_885012108020_4.7uF
*******
.subckt 1206_885012108021_10uF 1 2
Rser 1 3 0.00349318752029
Lser 2 4 6.43774867E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012108021_10uF
*******
.subckt 1210_885012109012_4.7uF 1 2
Rser 1 3 0.0033906445918
Lser 2 4 3.01326093E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012109012_4.7uF
*******
.subckt 1210_885012109013_10uF 1 2
Rser 1 3 0.00241697975791
Lser 2 4 8.77086276E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1210_885012109013_10uF
*******
.subckt 1210_885012109014_22uF 1 2
Rser 1 3 0.00268514753558
Lser 2 4 9.0689132E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1210_885012109014_22uF
*******
.subckt 1210_885012109015_22uF 1 2
Rser 1 3 0.00734474129923
Lser 2 4 1.236549611E-09
C1 3 4 0.000022
Rpar 3 4 5000000
.ends 1210_885012109015_22uF
*******
.subckt 0402_885012205038_100pF 1 2
Rser 1 3 0.81685
Lser 2 4 0.00000000015556
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012205038_100pF
*******
.subckt 0402_885012205039_150pF 1 2
Rser 1 3 0.63099
Lser 2 4 0.00000000012911
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012205039_150pF
*******
.subckt 0402_885012205040_220pF 1 2
Rser 1 3 0.56531
Lser 2 4 0.00000000019063
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012205040_220pF
*******
.subckt 0402_885012205041_330pF 1 2
Rser 1 3 0.47337
Lser 2 4 0.00000000018072
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012205041_330pF
*******
.subckt 0402_885012205042_470pF 1 2
Rser 1 3 0.34662
Lser 2 4 0.00000000017045
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012205042_470pF
*******
.subckt 0402_885012205043_680pF 1 2
Rser 1 3 0.26546
Lser 2 4 0.00000000014081
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0402_885012205043_680pF
*******
.subckt 0402_885012205044_1nF 1 2
Rser 1 3 0.2145
Lser 2 4 0.000000000153
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205044_1nF
*******
.subckt 0402_885012205045_1.5nF 1 2
Rser 1 3 0.20285
Lser 2 4 0.00000000025723
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0402_885012205045_1.5nF
*******
.subckt 0402_885012205046_2.2nF 1 2
Rser 1 3 0.16081
Lser 2 4 0.00000000018799
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0402_885012205046_2.2nF
*******
.subckt 0402_885012205047_3.3nF 1 2
Rser 1 3 0.12518
Lser 2 4 0.00000000020592
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0402_885012205047_3.3nF
*******
.subckt 0402_885012205048_4.7nF 1 2
Rser 1 3 0.09048
Lser 2 4 0.00000000014994
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205048_4.7nF
*******
.subckt 0402_885012205049_6.8nF 1 2
Rser 1 3 0.071
Lser 2 4 0.00000000019016
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0402_885012205049_6.8nF
*******
.subckt 0402_885012205050_10nF 1 2
Rser 1 3 0.0592
Lser 2 4 0.00000000014515
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0402_885012205050_10nF
*******
.subckt 0402_885012205051_15nF 1 2
Rser 1 3 0.03784
Lser 2 4 0.00000000020335
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0402_885012205051_15nF
*******
.subckt 0402_885012205052_22nF 1 2
Rser 1 3 0.0548
Lser 2 4 0.00000000019383
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0402_885012205052_22nF
*******
.subckt 0402_885012205053_33nF 1 2
Rser 1 3 0.03148
Lser 2 4 0.0000000002517
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0402_885012205053_33nF
*******
.subckt 0402_885012205054_47nF 1 2
Rser 1 3 0.02098
Lser 2 4 0.00000000019891
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0402_885012205054_47nF
*******
.subckt 0402_885012205085_100nF 1 2
Rser 1 3 0.035
Lser 2 4 7.65573672E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205085_100nF
*******
.subckt 0402_885012205085R_100nF 1 2
Rser 1 3 0.035
Lser 2 4 7.65573672E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205085R_100nF
*******
.subckt 0603_885012206053_100pF 1 2
Rser 1 3 0.91003
Lser 2 4 0.00000000024509
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206053_100pF
*******
.subckt 0603_885012206054_150pF 1 2
Rser 1 3 0.68385
Lser 2 4 0.00000000029018
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012206054_150pF
*******
.subckt 0603_885012206055_220pF 1 2
Rser 1 3 0.58631
Lser 2 4 0.00000000033037
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012206055_220pF
*******
.subckt 0603_885012206056_330pF 1 2
Rser 1 3 0.42401
Lser 2 4 0.00000000033129
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206056_330pF
*******
.subckt 0603_885012206057_470pF 1 2
Rser 1 3 0.34594
Lser 2 4 0.00000000033084
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206057_470pF
*******
.subckt 0603_885012206058_680pF 1 2
Rser 1 3 0.29796
Lser 2 4 0.00000000037378
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206058_680pF
*******
.subckt 0603_885012206059_1nF 1 2
Rser 1 3 0.22136
Lser 2 4 0.00000000036253
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206059_1nF
*******
.subckt 0603_885012206060_1.5nF 1 2
Rser 1 3 0.18842
Lser 2 4 0.00000000033832
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206060_1.5nF
*******
.subckt 0603_885012206061_2.2nF 1 2
Rser 1 3 0.12731
Lser 2 4 0.00000000032293
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012206061_2.2nF
*******
.subckt 0603_885012206062_3.3nF 1 2
Rser 1 3 0.09865
Lser 2 4 0.0000000003316
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206062_3.3nF
*******
.subckt 0603_885012206063_4.7nF 1 2
Rser 1 3 0.08147
Lser 2 4 0.0000000002893
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206063_4.7nF
*******
.subckt 0603_885012206064_6.8nF 1 2
Rser 1 3 0.08487
Lser 2 4 0.00000000036849
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206064_6.8nF
*******
.subckt 0603_885012206065_10nF 1 2
Rser 1 3 0.05893
Lser 2 4 0.00000000037916
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206065_10nF
*******
.subckt 0603_885012206066_15nF 1 2
Rser 1 3 0.0473
Lser 2 4 0.00000000030093
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0603_885012206066_15nF
*******
.subckt 0603_885012206067_22nF 1 2
Rser 1 3 0.03101
Lser 2 4 0.00000000028048
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885012206067_22nF
*******
.subckt 0603_885012206068_33nF 1 2
Rser 1 3 0.0232
Lser 2 4 0.00000000033089
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0603_885012206068_33nF
*******
.subckt 0603_885012206069_47nF 1 2
Rser 1 3 0.01832
Lser 2 4 0.0000000002418
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0603_885012206069_47nF
*******
.subckt 0603_885012206070_68nF 1 2
Rser 1 3 0.01712
Lser 2 4 0.00000000030682
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0603_885012206070_68nF
*******
.subckt 0603_885012206071_100nF 1 2
Rser 1 3 0.025
Lser 2 4 0.0000000008
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206071_100nF
*******
.subckt 0603_885012206071R_100nF 1 2
Rser 1 3 0.0189365521551
Lser 2 4 4.42668552E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206071R_100nF
*******
.subckt 0603_885012206072_150nF 1 2
Rser 1 3 0.0149181934238
Lser 2 4 3.31198563E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0603_885012206072_150nF
*******
.subckt 0603_885012206073_220nF 1 2
Rser 1 3 0.0109800094243
Lser 2 4 4.08100466E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012206073_220nF
*******
.subckt 0603_885012206074_330nF 1 2
Rser 1 3 0.0118150527569
Lser 2 4 4.48623546E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012206074_330nF
*******
.subckt 0603_885012206075_470nF 1 2
Rser 1 3 0.0100816359349
Lser 2 4 4.14055319E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012206075_470nF
*******
.subckt 0603_885012206075R_470nF 1 2
Rser 1 3 0.0100816359349
Lser 2 4 4.14055319E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012206075R_470nF
*******
.subckt 0603_885012206076_1uF 1 2
Rser 1 3 0.0073448307676
Lser 2 4 4.75503387E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0603_885012206076_1uF
*******
.subckt 0805_885012207054_100pF 1 2
Rser 1 3 0.90625
Lser 2 4 0.00000000029357
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207054_100pF
*******
.subckt 0805_885012207055_150pF 1 2
Rser 1 3 0.70433
Lser 2 4 0.00000000030352
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012207055_150pF
*******
.subckt 0805_885012207056_220pF 1 2
Rser 1 3 0.48805
Lser 2 4 0.00000000027764
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012207056_220pF
*******
.subckt 0805_885012207057_330pF 1 2
Rser 1 3 0.44753
Lser 2 4 0.00000000032997
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012207057_330pF
*******
.subckt 0805_885012207058_470pF 1 2
Rser 1 3 0.32032
Lser 2 4 0.0000000002982
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207058_470pF
*******
.subckt 0805_885012207059_680pF 1 2
Rser 1 3 0.25951
Lser 2 4 0.00000000036777
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012207059_680pF
*******
.subckt 0805_885012207060_1nF 1 2
Rser 1 3 0.20128
Lser 2 4 0.00000000029022
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207060_1nF
*******
.subckt 0805_885012207061_1.5nF 1 2
Rser 1 3 0.15833
Lser 2 4 0.00000000037277
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207061_1.5nF
*******
.subckt 0805_885012207062_2.2nF 1 2
Rser 1 3 0.11878
Lser 2 4 0.00000000036877
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012207062_2.2nF
*******
.subckt 0805_885012207063_3.3nF 1 2
Rser 1 3 0.10404
Lser 2 4 0.00000000034071
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207063_3.3nF
*******
.subckt 0805_885012207064_4.7nF 1 2
Rser 1 3 0.07475
Lser 2 4 0.00000000024317
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012207064_4.7nF
*******
.subckt 0805_885012207065_6.8nF 1 2
Rser 1 3 0.08276
Lser 2 4 0.00000000032015
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0805_885012207065_6.8nF
*******
.subckt 0805_885012207066_10nF 1 2
Rser 1 3 0.06408
Lser 2 4 0.0000000002943
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207066_10nF
*******
.subckt 0805_885012207067_15nF 1 2
Rser 1 3 0.05208
Lser 2 4 0.00000000031399
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0805_885012207067_15nF
*******
.subckt 0805_885012207068_22nF 1 2
Rser 1 3 0.0486328028818
Lser 2 4 0.00000000041
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0805_885012207068_22nF
*******
.subckt 0805_885012207069_33nF 1 2
Rser 1 3 0.0330484373884
Lser 2 4 0.00000000041
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0805_885012207069_33nF
*******
.subckt 0805_885012207070_47nF 1 2
Rser 1 3 0.0298909488495
Lser 2 4 0.00000000038
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0805_885012207070_47nF
*******
.subckt 0805_885012207071_68nF 1 2
Rser 1 3 0.0247
Lser 2 4 0.00000000027034
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0805_885012207071_68nF
*******
.subckt 0805_885012207072_100nF 1 2
Rser 1 3 0.0172819633028
Lser 2 4 0.00000000035
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207072_100nF
*******
.subckt 0805_885012207073_150nF 1 2
Rser 1 3 0.0145783171748
Lser 2 4 0.00000000035
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0805_885012207073_150nF
*******
.subckt 0805_885012207074_220nF 1 2
Rser 1 3 0.0111697818844
Lser 2 4 0.00000000042
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885012207074_220nF
*******
.subckt 0805_885012207075_330nF 1 2
Rser 1 3 0.00939488017121
Lser 2 4 0.000000000283
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885012207075_330nF
*******
.subckt 0805_885012207076_470nF 1 2
Rser 1 3 0.00781019032257
Lser 2 4 0.00000000049
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0805_885012207076_470nF
*******
.subckt 0805_885012207077_680nF 1 2
Rser 1 3 0.00783503615977
Lser 2 4 0.00000000053
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0805_885012207077_680nF
*******
.subckt 0805_885012207078_1uF 1 2
Rser 1 3 0.00804838198988
Lser 2 4 2.69843792E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885012207078_1uF
*******
.subckt 0805_885012207079_2.2uF 1 2
Rser 1 3 0.00468718250549
Lser 2 4 2.80891331E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012207079_2.2uF
*******
.subckt 1206_885012208042_220pF 1 2
Rser 1 3 0.58352
Lser 2 4 0.00000000032083
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012208042_220pF
*******
.subckt 1206_885012208043_330pF 1 2
Rser 1 3 0.50009
Lser 2 4 0.00000000035086
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012208043_330pF
*******
.subckt 1206_885012208044_470pF 1 2
Rser 1 3 0.35551
Lser 2 4 0.0000000004724
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208044_470pF
*******
.subckt 1206_885012208045_680pF 1 2
Rser 1 3 0.32598
Lser 2 4 0.0000000006527
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012208045_680pF
*******
.subckt 1206_885012208046_1nF 1 2
Rser 1 3 0.23112
Lser 2 4 0.00000000050124
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208046_1nF
*******
.subckt 1206_885012208047_1.5nF 1 2
Rser 1 3 0.17032
Lser 2 4 0.00000000040983
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012208047_1.5nF
*******
.subckt 1206_885012208048_2.2nF 1 2
Rser 1 3 0.11761
Lser 2 4 0.00000000058541
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012208048_2.2nF
*******
.subckt 1206_885012208049_3.3nF 1 2
Rser 1 3 0.12683
Lser 2 4 0.00000000044431
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012208049_3.3nF
*******
.subckt 1206_885012208050_4.7nF 1 2
Rser 1 3 0.07742
Lser 2 4 0.00000000042481
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208050_4.7nF
*******
.subckt 1206_885012208051_6.8nF 1 2
Rser 1 3 0.0893088703811
Lser 2 4 5.44959228E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012208051_6.8nF
*******
.subckt 1206_885012208052_10nF 1 2
Rser 1 3 0.355515780687
Lser 2 4 4.90239917E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208052_10nF
*******
.subckt 1206_885012208053_15nF 1 2
Rser 1 3 0.05086
Lser 2 4 0.00000000064474
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1206_885012208053_15nF
*******
.subckt 1206_885012208054_22nF 1 2
Rser 1 3 0.04388
Lser 2 4 0.00000000043595
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1206_885012208054_22nF
*******
.subckt 1206_885012208055_33nF 1 2
Rser 1 3 0.05974
Lser 2 4 0.00000000046935
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1206_885012208055_33nF
*******
.subckt 1206_885012208056_47nF 1 2
Rser 1 3 0.05553
Lser 2 4 0.00000000049393
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1206_885012208056_47nF
*******
.subckt 1206_885012208057_68nF 1 2
Rser 1 3 0.03879
Lser 2 4 0.00000000044546
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 1206_885012208057_68nF
*******
.subckt 1206_885012208058_100nF 1 2
Rser 1 3 0.0232208356231
Lser 2 4 5.59299026E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885012208058_100nF
*******
.subckt 1206_885012208059_150nF 1 2
Rser 1 3 0.0179362383614
Lser 2 4 5.89126458E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1206_885012208059_150nF
*******
.subckt 1206_885012208060_220nF 1 2
Rser 1 3 0.0124482582844
Lser 2 4 5.568771E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1206_885012208060_220nF
*******
.subckt 1206_885012208061_330nF 1 2
Rser 1 3 0.0123070322618
Lser 2 4 7.16267872E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1206_885012208061_330nF
*******
.subckt 1206_885012208062_470nF 1 2
Rser 1 3 0.0100846165597
Lser 2 4 7.45549291E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1206_885012208062_470nF
*******
.subckt 1206_885012208063_680nF 1 2
Rser 1 3 0.00806863562842
Lser 2 4 7.09595993E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1206_885012208063_680nF
*******
.subckt 1206_885012208064_1uF 1 2
Rser 1 3 0.00633398843665
Lser 2 4 7.50258152E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885012208064_1uF
*******
.subckt 1206_885012208065_1.5uF 1 2
Rser 1 3 0.00655648262409
Lser 2 4 8.57454998E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 1206_885012208065_1.5uF
*******
.subckt 1206_885012208066_2.2uF 1 2
Rser 1 3 0.00520440828302
Lser 2 4 7.87876644E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012208066_2.2uF
*******
.subckt 1206_885012208067_3.3uF 1 2
Rser 1 3 0.00537091922132
Lser 2 4 8.20379233E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012208067_3.3uF
*******
.subckt 1206_885012208068_4.7uF 1 2
Rser 1 3 0.00336451412099
Lser 2 4 7.97503693E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1206_885012208068_4.7uF
*******
.subckt 1206_885012208069_10uF 1 2
Rser 1 3 0.0039007012861
Lser 2 4 0.00000000055
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012208069_10uF
*******
.subckt 1210_885012209015_1nF 1 2
Rser 1 3 0.23064
Lser 2 4 0.00000000009004
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885012209015_1nF
*******
.subckt 1210_885012209016_2.2nF 1 2
Rser 1 3 0.15
Lser 2 4 0.0000000009
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1210_885012209016_2.2nF
*******
.subckt 1210_885012209017_10nF 1 2
Rser 1 3 0.07411
Lser 2 4 0.00000000018051
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1210_885012209017_10nF
*******
.subckt 1210_885012209018_22nF 1 2
Rser 1 3 0.06131
Lser 2 4 0.00000000020837
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1210_885012209018_22nF
*******
.subckt 1210_885012209019_100nF 1 2
Rser 1 3 0.0209574310072
Lser 2 4 5.49171232E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1210_885012209019_100nF
*******
.subckt 1210_885012209020_220nF 1 2
Rser 1 3 0.0109918196754
Lser 2 4 5.14177759E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1210_885012209020_220nF
*******
.subckt 1210_885012209021_330nF 1 2
Rser 1 3 0.00972375707294
Lser 2 4 5.4771949E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1210_885012209021_330nF
*******
.subckt 1210_885012209022_470nF 1 2
Rser 1 3 0.00740093895541
Lser 2 4 5.16300103E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1210_885012209022_470nF
*******
.subckt 1210_885012209023_680nF 1 2
Rser 1 3 0.00560873026626
Lser 2 4 5.62947674E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1210_885012209023_680nF
*******
.subckt 1210_885012209024_1uF 1 2
Rser 1 3 0.00434521559376
Lser 2 4 3.4952573E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209024_1uF
*******
.subckt 1210_885012209025_2.2uF 1 2
Rser 1 3 0.003755566195
Lser 2 4 4.76192409E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1210_885012209025_2.2uF
*******
.subckt 1210_885012209026_3.3uF 1 2
Rser 1 3 0.0037725139254
Lser 2 4 4.43584901E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1210_885012209026_3.3uF
*******
.subckt 1210_885012209027_4.7uF 1 2
Rser 1 3 0.00334303070776
Lser 2 4 4.2432524E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012209027_4.7uF
*******
.subckt 1210_885012209028_10uF 1 2
Rser 1 3 0.0026086390311
Lser 2 4 8.94000611E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1210_885012209028_10uF
*******
.subckt 1210_885012209074_22uF 1 2
Rser 1 3 0.0043
Lser 2 4 0.000000001
C1 3 4 0.000022
Rpar 3 4 5000000
.ends 1210_885012209074_22uF
*******
.subckt 1812_885012210005_4.7nF 1 2
Rser 1 3 0.0828
Lser 2 4 0.00000000018862
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1812_885012210005_4.7nF
*******
.subckt 1812_885012210006_10nF 1 2
Rser 1 3 0.07693
Lser 2 4 0.00000000053548
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012210006_10nF
*******
.subckt 1812_885012210007_47nF 1 2
Rser 1 3 0.03468
Lser 2 4 0.00000000076842
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1812_885012210007_47nF
*******
.subckt 1812_885012210008_100nF 1 2
Rser 1 3 0.037008688888
Lser 2 4 6.73793576E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1812_885012210008_100nF
*******
.subckt 1812_885012210009_330nF 1 2
Rser 1 3 0.01427157177
Lser 2 4 4.80558989E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1812_885012210009_330nF
*******
.subckt 1812_885012210010_470nF 1 2
Rser 1 3 0.00985565119595
Lser 2 4 4.00753105E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1812_885012210010_470nF
*******
.subckt 1812_885012210011_680nF 1 2
Rser 1 3 0.00784524987635
Lser 2 4 4.30816782E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1812_885012210011_680nF
*******
.subckt 1812_885012210012_1uF 1 2
Rser 1 3 0.014
Lser 2 4 0.000000001
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1812_885012210012_1uF
*******
.subckt 0201_885012004001_100pF 1 2
Rser 1 3 0.2125
Lser 2 4 0.00000000025
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0201_885012004001_100pF
*******
.subckt 0201_885012204004_10nF 1 2
Rser 1 3 0.0709
Lser 2 4 0.00000000018
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012204004_10nF
*******
.subckt 0201_885012104005_100nF 1 2
Rser 1 3 0.0287
Lser 2 4 0.00000000015
C1 3 4 0.0000001
Rpar 3 4 500000000
.ends 0201_885012104005_100nF
*******
.subckt 0201_885012104008_4.7nF 1 2
Rser 1 3 0.093
Lser 2 4 0.000000000212
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0201_885012104008_4.7nF
*******
.subckt 0201_885012004003_1.5pF 1 2
Rser 1 3 0.8126
Lser 2 4 0.00000000022
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0201_885012004003_1.5pF
*******
.subckt 0201_885012004004_10pF 1 2
Rser 1 3 0.6361
Lser 2 4 0.00000000022
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0201_885012004004_10pF
*******
.subckt 0201_885012004005_12pF 1 2
Rser 1 3 0.4731
Lser 2 4 0.00000000021
C1 3 4 0.000000000012
Rpar 3 4 10000000000
.ends 0201_885012004005_12pF
*******
.subckt 0201_885012004006_15pF 1 2
Rser 1 3 0.4471
Lser 2 4 0.00000000025
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0201_885012004006_15pF
*******
.subckt 0201_885012004007_18pF 1 2
Rser 1 3 0.4894
Lser 2 4 0.000000000295
C1 3 4 0.000000000018
Rpar 3 4 10000000000
.ends 0201_885012004007_18pF
*******
.subckt 0201_885012004008_22pF 1 2
Rser 1 3 0.5288
Lser 2 4 0.00000000026
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0201_885012004008_22pF
*******
.subckt 0201_885012004009_33pF 1 2
Rser 1 3 0.3381
Lser 2 4 0.000000000257
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0201_885012004009_33pF
*******
.subckt 0201_885012004010_47pF 1 2
Rser 1 3 0.241
Lser 2 4 0.0000000002
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0201_885012004010_47pF
*******
.subckt 0201_885012204006_1nF 1 2
Rser 1 3 0.2367
Lser 2 4 0.000000000173
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0201_885012204006_1nF
*******
.subckt 0201_885012104014_10nF 1 2
Rser 1 3 0.0639
Lser 2 4 0.00000000021
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012104014_10nF
*******
.subckt 2220_885012214004_10uF 1 2
Rser 1 3 0.003
Lser 2 4 0.0000000012
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 2220_885012214004_10uF
*******
.subckt 0603_885012106030_1uF 1 2
Rser 1 3 0.013
Lser 2 4 0.0000000008
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0603_885012106030_1uF
*******
.subckt 0402_885012005007_10pF 1 2
Rser 1 3 0.494547705824
Lser 2 4 3.67389142E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005007_10pF
*******
.subckt 0402_885012005008_15pF 1 2
Rser 1 3 0.388190780491
Lser 2 4 3.17307789E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885012005008_15pF
*******
.subckt 0402_885012005009_22pF 1 2
Rser 1 3 0.316230222598
Lser 2 4 2.88077478E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885012005009_22pF
*******
.subckt 0402_885012005010_33pF 1 2
Rser 1 3 0.249324470259
Lser 2 4 2.84730223E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005010_33pF
*******
.subckt 0402_885012005011_47pF 1 2
Rser 1 3 0.235686289563
Lser 2 4 2.78272514E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005011_47pF
*******
.subckt 0402_885012005012_68pF 1 2
Rser 1 3 0.188011183755
Lser 2 4 2.62979806E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005012_68pF
*******
.subckt 0402_885012005013_100pF 1 2
Rser 1 3 0.145490051878
Lser 2 4 2.5124412E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005013_100pF
*******
.subckt 0402_885012005014_150pF 1 2
Rser 1 3 0.102893245885
Lser 2 4 2.1894381E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012005014_150pF
*******
.subckt 0402_885012005015_220pF 1 2
Rser 1 3 0.0932691679838
Lser 2 4 1.50271806E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012005015_220pF
*******
.subckt 0402_885012005016_330pF 1 2
Rser 1 3 0.0893241489871
Lser 2 4 3.29295953E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012005016_330pF
*******
.subckt 0402_885012005017_470pF 1 2
Rser 1 3 0.0149178531097
Lser 2 4 3.26241368E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012005017_470pF
*******
.subckt 0402_885012005018_1nF 1 2
Rser 1 3 0.0157004412396
Lser 2 4 3.37941862E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012005018_1nF
*******
.subckt 0603_885012006001_4.7pF 1 2
Rser 1 3 0.307143942354
Lser 2 4 3.18870536E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0603_885012006001_4.7pF
*******
.subckt 0603_885012006002_10pF 1 2
Rser 1 3 0.668
Lser 2 4 0.00000000056
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006002_10pF
*******
.subckt 0603_885012006003_15pF 1 2
Rser 1 3 0.318625808147
Lser 2 4 7.07424269E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006003_15pF
*******
.subckt 0603_885012006004_22pF 1 2
Rser 1 3 0.34819611654
Lser 2 4 7.75018519E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006004_22pF
*******
.subckt 0603_885012006005_33pF 1 2
Rser 1 3 0.266845513997
Lser 2 4 8.03723788E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006005_33pF
*******
.subckt 0603_885012006006_47pF 1 2
Rser 1 3 0.196782783005
Lser 2 4 7.59426691E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006006_47pF
*******
.subckt 0603_885012006007_68pF 1 2
Rser 1 3 0.153641735222
Lser 2 4 7.22489136E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006007_68pF
*******
.subckt 0603_885012006008_100pF 1 2
Rser 1 3 0.110129832129
Lser 2 4 6.73785263E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006008_100pF
*******
.subckt 0603_885012006009_150pF 1 2
Rser 1 3 0.0793891689318
Lser 2 4 6.22415559E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006009_150pF
*******
.subckt 0603_885012006010_220pF 1 2
Rser 1 3 0.088220302088
Lser 2 4 6.95492511E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012006010_220pF
*******
.subckt 0603_885012006011_330pF 1 2
Rser 1 3 0.0993151086205
Lser 2 4 4.18653134E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006011_330pF
*******
.subckt 0603_885012006012_470pF 1 2
Rser 1 3 0.0757443435992
Lser 2 4 3.66481782E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006012_470pF
*******
.subckt 0603_885012006013_680pF 1 2
Rser 1 3 0.0602766942369
Lser 2 4 3.26882078E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006013_680pF
*******
.subckt 0603_885012006014_1nF 1 2
Rser 1 3 0.0434067925003
Lser 2 4 4.09321859E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006014_1nF
*******
.subckt 0603_885012006015_2.2nF 1 2
Rser 1 3 0.0307077888885
Lser 2 4 3.39702907E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012006015_2.2nF
*******
.subckt 0603_885012006016_3.3nF 1 2
Rser 1 3 0.0275317919224
Lser 2 4 3.37901927E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012006016_3.3nF
*******
.subckt 0805_885012007001_15pF 1 2
Rser 1 3 0.322686614764
Lser 2 4 5.17792028E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007001_15pF
*******
.subckt 0805_885012007002_22pF 1 2
Rser 1 3 0.304017782882
Lser 2 4 6.06807592E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0805_885012007002_22pF
*******
.subckt 0805_885012007003_33pF 1 2
Rser 1 3 0.278413141435
Lser 2 4 5.73322702E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007003_33pF
*******
.subckt 0805_885012007004_100pF 1 2
Rser 1 3 0.144376756
Lser 2 4 4.19735168E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007004_100pF
*******
.subckt 0805_885012007005_150pF 1 2
Rser 1 3 0.132070069125
Lser 2 4 4.14007712E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007005_150pF
*******
.subckt 0805_885012007006_330pF 1 2
Rser 1 3 0.0858219234392
Lser 2 4 4.4258651E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007006_330pF
*******
.subckt 0805_885012007007_470pF 1 2
Rser 1 3 0.0754569114616
Lser 2 4 4.35286885E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007007_470pF
*******
.subckt 0805_885012007008_1nF 1 2
Rser 1 3 0.0525130505561
Lser 2 4 4.16381481E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007008_1nF
*******
.subckt 0805_885012007009_10nF 1 2
Rser 1 3 0.0143302506767
Lser 2 4 2.53788056E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012007009_10nF
*******
.subckt 1206_885012008001_10pF 1 2
Rser 1 3 0.446014275484
Lser 2 4 5.73571915E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1206_885012008001_10pF
*******
.subckt 1206_885012008002_22pF 1 2
Rser 1 3 0.299003095867
Lser 2 4 5.45254376E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1206_885012008002_22pF
*******
.subckt 1206_885012008003_47pF 1 2
Rser 1 3 0.21040740508
Lser 2 4 5.6609278E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885012008003_47pF
*******
.subckt 1206_885012008004_100pF 1 2
Rser 1 3 0.167865253643
Lser 2 4 4.85486348E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008004_100pF
*******
.subckt 1206_885012008005_470pF 1 2
Rser 1 3 0.115247377385
Lser 2 4 4.7229295E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012008005_470pF
*******
.subckt 1206_885012008006_2.2nF 1 2
Rser 1 3 0.0350339469969
Lser 2 4 1.042313537E-12
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012008006_2.2nF
*******
.subckt 1206_885012008007_6.8nF 1 2
Rser 1 3 0.0298615638448
Lser 2 4 9.14635803E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008007_6.8nF
*******
.subckt 1206_885012008008_10nF 1 2
Rser 1 3 0.0249778783357
Lser 2 4 9.13131263E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008008_10nF
*******
.subckt 1206_885012008009_22nF 1 2
Rser 1 3 0.011442234975
Lser 2 4 8.6240711E-10
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1206_885012008009_22nF
*******
.subckt 1206_885012008010_33nF 1 2
Rser 1 3 0.0092860021616
Lser 2 4 8.63894198E-10
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1206_885012008010_33nF
*******
.subckt 0402_885012105009_68nF 1 2
Rser 1 3 0.0638704519417
Lser 2 4 2.20630867E-10
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0402_885012105009_68nF
*******
.subckt 0402_885012105010_100nF 1 2
Rser 1 3 0.0268043216773
Lser 2 4 3.11178988E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012105010_100nF
*******
.subckt 0402_885012105011_220nF 1 2
Rser 1 3 0.0122717751401
Lser 2 4 3.48439745E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0402_885012105011_220nF
*******
.subckt 0402_885012105012_1uF 1 2
Rser 1 3 0.00986403339919
Lser 2 4 3.2821055E-10
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0402_885012105012_1uF
*******
.subckt 0402_885012105013_2.2uF 1 2
Rser 1 3 0.009771521005
Lser 2 4 3.03733414E-10
C1 3 4 0.0000022
Rpar 3 4 20000000
.ends 0402_885012105013_2.2uF
*******
.subckt 0603_885012106007_330nF 1 2
Rser 1 3 0.0111038975002
Lser 2 4 3.20933284E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012106007_330nF
*******
.subckt 0603_885012106008_470nF 1 2
Rser 1 3 0.00949633292517
Lser 2 4 2.70539302E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0603_885012106008_470nF
*******
.subckt 0603_885012106009_680nF 1 2
Rser 1 3 0.0112015362567
Lser 2 4 3.50610132E-10
C1 3 4 0.00000068
Rpar 3 4 200000000
.ends 0603_885012106009_680nF
*******
.subckt 0603_885012106010_1uF 1 2
Rser 1 3 0.00802031801588
Lser 2 4 3.00240209E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012106010_1uF
*******
.subckt 0603_885012106011_2.2uF 1 2
Rser 1 3 0.00618507884481
Lser 2 4 2.53136283E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0603_885012106011_2.2uF
*******
.subckt 0603_885012106012_4.7uF 1 2
Rser 1 3 0.00455496693599
Lser 2 4 5.03384516E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0603_885012106012_4.7uF
*******
.subckt 0805_885012107007_2.2uF 1 2
Rser 1 3 0.00451361812717
Lser 2 4 2.56807852E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012107007_2.2uF
*******
.subckt 0805_885012107008_3.3uF 1 2
Rser 1 3 0.00416445411098
Lser 2 4 3.00167169E-10
C1 3 4 0.0000033
Rpar 3 4 30000000
.ends 0805_885012107008_3.3uF
*******
.subckt 0805_885012107009_4.7uF 1 2
Rser 1 3 0.00333037459922
Lser 2 4 2.41667028E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0805_885012107009_4.7uF
*******
.subckt 0805_885012107010_10uF 1 2
Rser 1 3 0.00257315295813
Lser 2 4 4.16651033E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 0805_885012107010_10uF
*******
.subckt 0805_885012107011_22uF 1 2
Rser 1 3 0.00309713657007
Lser 2 4 2.86347556E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 0805_885012107011_22uF
*******
.subckt 1206_885012108006_2.2uF 1 2
Rser 1 3 0.00715208568262
Lser 2 4 5.64041345E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012108006_2.2uF
*******
.subckt 1206_885012108007_3.3uF 1 2
Rser 1 3 0.00529476260464
Lser 2 4 6.12367847E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012108007_3.3uF
*******
.subckt 1206_885012108008_4.7uF 1 2
Rser 1 3 0.00610205096672
Lser 2 4 5.17669274E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012108008_4.7uF
*******
.subckt 1206_885012108009_6.8uF 1 2
Rser 1 3 0.00416216687199
Lser 2 4 6.95534046E-10
C1 3 4 0.0000068
Rpar 3 4 20000000
.ends 1206_885012108009_6.8uF
*******
.subckt 1206_885012108010_10uF 1 2
Rser 1 3 0.00362327531378
Lser 2 4 0.0000000008
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1206_885012108010_10uF
*******
.subckt 1206_885012108011_22uF 1 2
Rser 1 3 0.00240452659004
Lser 2 4 8.37875791E-10
C1 3 4 0.000022
Rpar 3 4 5000000
.ends 1206_885012108011_22uF
*******
.subckt 1206_885012108012_47uF 1 2
Rser 1 3 0.0027428064885
Lser 2 4 0.0000000008
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1206_885012108012_47uF
*******
.subckt 1210_885012109005_10uF 1 2
Rser 1 3 0.00250479636867
Lser 2 4 7.49918881E-10
C1 3 4 0.00001
Rpar 3 4 50000000
.ends 1210_885012109005_10uF
*******
.subckt 1210_885012109006_22uF 1 2
Rser 1 3 0.00272955719838
Lser 2 4 9.31961125E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1210_885012109006_22uF
*******
.subckt 1210_885012109007_47uF 1 2
Rser 1 3 0.00210105515092
Lser 2 4 0.0000000009
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1210_885012109007_47uF
*******
.subckt 0402_885012205001_100pF 1 2
Rser 1 3 0.78619
Lser 2 4 0.00000000015138
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012205001_100pF
*******
.subckt 0402_885012205002_220pF 1 2
Rser 1 3 0.5727
Lser 2 4 1.77695991E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012205002_220pF
*******
.subckt 0402_885012205003_330pF 1 2
Rser 1 3 0.43753
Lser 2 4 0.00000000020201
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012205003_330pF
*******
.subckt 0402_885012205004_470pF 1 2
Rser 1 3 0.33537
Lser 2 4 0.00000000018013
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012205004_470pF
*******
.subckt 0402_885012205005_680pF 1 2
Rser 1 3 0.26133
Lser 2 4 0.00000000015756
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0402_885012205005_680pF
*******
.subckt 0402_885012205006_1nF 1 2
Rser 1 3 0.19089
Lser 2 4 0.00000000017743
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205006_1nF
*******
.subckt 0402_885012205007_1.5nF 1 2
Rser 1 3 0.16721
Lser 2 4 0.00000000024076
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0402_885012205007_1.5nF
*******
.subckt 0402_885012205008_2.2nF 1 2
Rser 1 3 0.11524
Lser 2 4 0.000000000227222
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0402_885012205008_2.2nF
*******
.subckt 0402_885012205009_3.3nF 1 2
Rser 1 3 0.0897
Lser 2 4 0.00000000023518
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0402_885012205009_3.3nF
*******
.subckt 0402_885012205010_4.7nF 1 2
Rser 1 3 0.05632
Lser 2 4 0.00000000018931
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205010_4.7nF
*******
.subckt 0402_885012205011_6.8nF 1 2
Rser 1 3 0.04164
Lser 2 4 0.00000000021064
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0402_885012205011_6.8nF
*******
.subckt 0402_885012205012_10nF 1 2
Rser 1 3 0.0531398956639
Lser 2 4 0.00000000022
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0402_885012205012_10nF
*******
.subckt 0402_885012205013_15nF 1 2
Rser 1 3 0.03039
Lser 2 4 0.00000000022583
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0402_885012205013_15nF
*******
.subckt 0402_885012205014_22nF 1 2
Rser 1 3 0.01645
Lser 2 4 0.00000000020049
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0402_885012205014_22nF
*******
.subckt 0402_885012205015_33nF 1 2
Rser 1 3 0.00701
Lser 2 4 0.00000000023581
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0402_885012205015_33nF
*******
.subckt 0402_885012205016_47nF 1 2
Rser 1 3 0.0071
Lser 2 4 0.0000000002065
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0402_885012205016_47nF
*******
.subckt 0402_885012205017_68nF 1 2
Rser 1 3 0.01539
Lser 2 4 0.00000000023044
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0402_885012205017_68nF
*******
.subckt 0402_885012205018_100nF 1 2
Rser 1 3 0.0183525691398
Lser 2 4 3.07541467E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205018_100nF
*******
.subckt 0603_885012206003_100pF 1 2
Rser 1 3 0.86219
Lser 2 4 0.00000000020992
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206003_100pF
*******
.subckt 0603_885012206004_220pF 1 2
Rser 1 3 0.55667
Lser 2 4 0.00000000030069
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012206004_220pF
*******
.subckt 0603_885012206005_330pF 1 2
Rser 1 3 0.43756
Lser 2 4 0.00000000026062
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206005_330pF
*******
.subckt 0603_885012206006_470pF 1 2
Rser 1 3 0.37246
Lser 2 4 0.00000000030107
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206006_470pF
*******
.subckt 0603_885012206007_680pF 1 2
Rser 1 3 0.31851
Lser 2 4 0.00000000040239
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206007_680pF
*******
.subckt 0603_885012206008_1nF 1 2
Rser 1 3 0.24958
Lser 2 4 0.00000000040399
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206008_1nF
*******
.subckt 0603_885012206009_1.5nF 1 2
Rser 1 3 0.20086
Lser 2 4 0.00000000033824
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206009_1.5nF
*******
.subckt 0603_885012206010_2.2nF 1 2
Rser 1 3 0.14948
Lser 2 4 0.00000000033334
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012206010_2.2nF
*******
.subckt 0603_885012206011_3.3nF 1 2
Rser 1 3 0.12415
Lser 2 4 0.00000000032537
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206011_3.3nF
*******
.subckt 0603_885012206012_4.7nF 1 2
Rser 1 3 0.07518
Lser 2 4 0.0000000003009
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206012_4.7nF
*******
.subckt 0603_885012206013_6.8nF 1 2
Rser 1 3 0.07031
Lser 2 4 0.00000000039053
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206013_6.8nF
*******
.subckt 0603_885012206014_10nF 1 2
Rser 1 3 0.04641
Lser 2 4 0.00000000025735
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206014_10nF
*******
.subckt 0603_885012206015_15nF 1 2
Rser 1 3 0.03908
Lser 2 4 0.00000000026071
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0603_885012206015_15nF
*******
.subckt 0603_885012206016_22nF 1 2
Rser 1 3 0.02302
Lser 2 4 0.00000000023719
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885012206016_22nF
*******
.subckt 0603_885012206017_33nF 1 2
Rser 1 3 0.01243
Lser 2 4 0.00000000025982
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0603_885012206017_33nF
*******
.subckt 0603_885012206018_47nF 1 2
Rser 1 3 0.01343
Lser 2 4 0.00000000024476
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0603_885012206018_47nF
*******
.subckt 0603_885012206019_68nF 1 2
Rser 1 3 0.0155
Lser 2 4 0.00000000030737
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0603_885012206019_68nF
*******
.subckt 0603_885012206020_100nF 1 2
Rser 1 3 0.0188883213835
Lser 2 4 4.53593763E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206020_100nF
*******
.subckt 0603_885012206021_150nF 1 2
Rser 1 3 0.0221138242279
Lser 2 4 4.07625742E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0603_885012206021_150nF
*******
.subckt 0603_885012206022_220nF 1 2
Rser 1 3 0.0146862228843
Lser 2 4 4.43010481E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012206022_220nF
*******
.subckt 0603_885012206023_330nF 1 2
Rser 1 3 0.0113479919005
Lser 2 4 4.48567636E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012206023_330nF
*******
.subckt 0603_885012206024_470nF 1 2
Rser 1 3 0.00961049589993
Lser 2 4 4.09343651E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0603_885012206024_470nF
*******
.subckt 0603_885012206025_680nF 1 2
Rser 1 3 0.00730055384166
Lser 2 4 4.35162169E-10
C1 3 4 0.00000068
Rpar 3 4 200000000
.ends 0603_885012206025_680nF
*******
.subckt 0603_885012206026_1uF 1 2
Rser 1 3 0.00743560640346
Lser 2 4 2.29632839E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012206026_1uF
*******
.subckt 0603_885012206027_2.2uF 1 2
Rser 1 3 0.00844425861819
Lser 2 4 2.90335669E-10
C1 3 4 0.0000022
Rpar 3 4 20000000
.ends 0603_885012206027_2.2uF
*******
.subckt 0805_885012207004_100pF 1 2
Rser 1 3 0.88264
Lser 2 4 0.00000000031858
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207004_100pF
*******
.subckt 0805_885012207005_220pF 1 2
Rser 1 3 0.50995
Lser 2 4 0.00000000027274
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012207005_220pF
*******
.subckt 0805_885012207006_470pF 1 2
Rser 1 3 0.31274
Lser 2 4 0.00000000031898
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207006_470pF
*******
.subckt 0805_885012207007_1nF 1 2
Rser 1 3 0.1905
Lser 2 4 0.00000000028002
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207007_1nF
*******
.subckt 0805_885012207008_1.5nF 1 2
Rser 1 3 0.16519
Lser 2 4 0.00000000038865
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207008_1.5nF
*******
.subckt 0805_885012207009_2.2nF 1 2
Rser 1 3 0.02478
Lser 2 4 0.00000000027522
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012207009_2.2nF
*******
.subckt 0805_885012207010_3.3nF 1 2
Rser 1 3 0.02239
Lser 2 4 0.00000000023565
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207010_3.3nF
*******
.subckt 0805_885012207011_10nF 1 2
Rser 1 3 0.04883
Lser 2 4 0.00000000031494
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207011_10nF
*******
.subckt 0805_885012207012_15nF 1 2
Rser 1 3 0.0512
Lser 2 4 0.00000000030048
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0805_885012207012_15nF
*******
.subckt 0805_885012207013_22nF 1 2
Rser 1 3 0.03858
Lser 2 4 0.00000000031876
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0805_885012207013_22nF
*******
.subckt 0805_885012207014_33nF 1 2
Rser 1 3 0.03079
Lser 2 4 0.00000000030588
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0805_885012207014_33nF
*******
.subckt 0805_885012207015_47nF 1 2
Rser 1 3 0.02162
Lser 2 4 0.0000000002672
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0805_885012207015_47nF
*******
.subckt 0805_885012207016_100nF 1 2
Rser 1 3 0.0162501221785
Lser 2 4 0.000000000375
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207016_100nF
*******
.subckt 0805_885012207017_150nF 1 2
Rser 1 3 0.0143154309487
Lser 2 4 4.47033542E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0805_885012207017_150nF
*******
.subckt 0805_885012207018_220nF 1 2
Rser 1 3 0.0114343175461
Lser 2 4 4.37838091E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885012207018_220nF
*******
.subckt 0805_885012207019_330nF 1 2
Rser 1 3 0.0106449562538
Lser 2 4 4.87419012E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885012207019_330nF
*******
.subckt 0805_885012207020_470nF 1 2
Rser 1 3 0.00823353483639
Lser 2 4 4.7697612E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0805_885012207020_470nF
*******
.subckt 0805_885012207021_680nF 1 2
Rser 1 3 0.00756100048721
Lser 2 4 5.19694932E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0805_885012207021_680nF
*******
.subckt 0805_885012207022_1uF 1 2
Rser 1 3 0.00779960743902
Lser 2 4 2.50116995E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885012207022_1uF
*******
.subckt 0805_885012207023_1.5uF 1 2
Rser 1 3 0.00625640838813
Lser 2 4 3.16162321E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 0805_885012207023_1.5uF
*******
.subckt 0805_885012207024_2.2uF 1 2
Rser 1 3 0.00498465718149
Lser 2 4 2.58299749E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012207024_2.2uF
*******
.subckt 0805_885012207025_4.7uF 1 2
Rser 1 3 0.00550893409975
Lser 2 4 2.51361537E-10
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0805_885012207025_4.7uF
*******
.subckt 0805_885012207026_10uF 1 2
Rser 1 3 0.00369416302331
Lser 2 4 5.01488494E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0805_885012207026_10uF
*******
.subckt 1206_885012208004_330pF 1 2
Rser 1 3 0.46442
Lser 2 4 0.00000000041059
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012208004_330pF
*******
.subckt 1206_885012208005_470pF 1 2
Rser 1 3 0.38435
Lser 2 4 0.00000000043066
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208005_470pF
*******
.subckt 1206_885012208006_1nF 1 2
Rser 1 3 0.22561
Lser 2 4 0.00000000045042
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208006_1nF
*******
.subckt 1206_885012208007_4.7nF 1 2
Rser 1 3 0.13666
Lser 2 4 0.00000000045064
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208007_4.7nF
*******
.subckt 1206_885012208008_10nF 1 2
Rser 1 3 0.06965
Lser 2 4 0.00000000068939
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208008_10nF
*******
.subckt 1206_885012208009_100nF 1 2
Rser 1 3 0.0244803326156
Lser 2 4 6.58788173E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885012208009_100nF
*******
.subckt 1206_885012208010_330nF 1 2
Rser 1 3 0.0123317635994
Lser 2 4 6.03276395E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1206_885012208010_330nF
*******
.subckt 1206_885012208011_470nF 1 2
Rser 1 3 0.010415539685
Lser 2 4 7.51451536E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1206_885012208011_470nF
*******
.subckt 1206_885012208012_680nF 1 2
Rser 1 3 0.00703741199294
Lser 2 4 7.17949052E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1206_885012208012_680nF
*******
.subckt 1206_885012208013_1uF 1 2
Rser 1 3 0.00648320483926
Lser 2 4 5.4243262E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885012208013_1uF
*******
.subckt 1206_885012208014_1.5uF 1 2
Rser 1 3 0.00911925278109
Lser 2 4 6.57782928E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 1206_885012208014_1.5uF
*******
.subckt 1206_885012208015_2.2uF 1 2
Rser 1 3 0.00662951285801
Lser 2 4 5.30235159E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012208015_2.2uF
*******
.subckt 1206_885012208016_3.3uF 1 2
Rser 1 3 0.00509978680029
Lser 2 4 6.27645723E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012208016_3.3uF
*******
.subckt 1206_885012208017_4.7uF 1 2
Rser 1 3 0.00357416297194
Lser 2 4 4.72459357E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012208017_4.7uF
*******
.subckt 1206_885012208018_10uF 1 2
Rser 1 3 0.00288901435933
Lser 2 4 7.48356777E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1206_885012208018_10uF
*******
.subckt 1206_885012208019_22uF 1 2
Rser 1 3 0.00343100506851
Lser 2 4 5.00393923E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1206_885012208019_22uF
*******
.subckt 1210_885012209001_47nF 1 2
Rser 1 3 0.03203
Lser 2 4 0.00000000012248
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1210_885012209001_47nF
*******
.subckt 1210_885012209002_220nF 1 2
Rser 1 3 0.0108946736088
Lser 2 4 5.13453415E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1210_885012209002_220nF
*******
.subckt 1210_885012209003_1uF 1 2
Rser 1 3 0.00441457708348
Lser 2 4 3.73414796E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209003_1uF
*******
.subckt 1210_885012209004_4.7uF 1 2
Rser 1 3 0.0051217091228
Lser 2 4 5.20978006E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012209004_4.7uF
*******
.subckt 1210_885012209005_10uF 1 2
Rser 1 3 0.00237372157538
Lser 2 4 7.95583466E-10
C1 3 4 0.00001
Rpar 3 4 100000000
.ends 1210_885012209005_10uF
*******
.subckt 1210_885012209006_22uF 1 2
Rser 1 3 0.0039
Lser 2 4 1.129373051E-09
C1 3 4 0.000022
Rpar 3 4 10000000
.ends 1210_885012209006_22uF
*******
.subckt 0201_885012104002_100nF 1 2
Rser 1 3 0.02596
Lser 2 4 0.00000000018
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0201_885012104002_100nF
*******
.subckt 0201_885012104006_220nF 1 2
Rser 1 3 0.02291
Lser 2 4 0.00000000015
C1 3 4 0.00000022
Rpar 3 4 200000000
.ends 0201_885012104006_220nF
*******
.subckt 0201_885012204005_10nF 1 2
Rser 1 3 0.0631
Lser 2 4 0.000000000217
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012204005_10nF
*******
.subckt 0201_885012104012_10nF 1 2
Rser 1 3 0.0632
Lser 2 4 0.000000000213
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012104012_10nF
*******
.subckt 0201_885012104013_47nF 1 2
Rser 1 3 0.06035
Lser 2 4 0.00000000022
C1 3 4 0.000000047
Rpar 3 4 2000000000
.ends 0201_885012104013_47nF
*******

