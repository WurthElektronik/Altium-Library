**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  HV SMT Dual Powerchoke
* Matchcode:              WE-DPC 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 5030_7448841010_1u  1  2  3  4  PARAMS:
+  Cww=6.54p
+  Rp1=1666
+  Cp1=0.725p
+  Lp1=0.9u
+  Rp2=1666
+  Cp2=0.725p
+  Lp2=0.9u
+  RDC1=0.032
+  RDC2=0.032
+  K=0.964365076099295
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841015_1.5u  1  2  3  4  PARAMS:
+  Cww=6.98p
+  Rp1=3088
+  Cp1=0.917p
+  Lp1=1.818u
+  Rp2=3088
+  Cp2=0.917p
+  Lp2=1.818u
+  RDC1=0.048
+  RDC2=0.048
+  K=0.972967967955095
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841022_2.2u  1  2  3  4  PARAMS:
+  Cww=7.46p
+  Rp1=4172
+  Cp1=1.291p
+  Lp1=2.312u
+  Rp2=4172
+  Cp2=1.291p
+  Lp2=2.312u
+  RDC1=0.05
+  RDC2=0.05
+  K=0.971175482691886
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841033_3.3u  1  2  3  4  PARAMS:
+  Cww=9.17p
+  Rp1=5673
+  Cp1=3.09p
+  Lp1=3.682u
+  Rp2=5673
+  Cp2=3.09p
+  Lp2=3.682u
+  RDC1=0.084
+  RDC2=0.084
+  K=0.980105127323626
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841047_4.7u  1  2  3  4  PARAMS:
+  Cww=10.01p
+  Rp1=7766
+  Cp1=2.824p
+  Lp1=5.957u
+  Rp2=7766
+  Cp2=2.824p
+  Lp2=5.957u
+  RDC1=0.102
+  RDC2=0.102
+  K=0.982831341995416
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841068_6.8u  1  2  3  4  PARAMS:
+  Cww=12.45p
+  Rp1=10491
+  Cp1=3.221p
+  Lp1=7.657u
+  Rp2=10491
+  Cp2=3.221p
+  Lp2=7.657u
+  RDC1=0.168
+  RDC2=0.168
+  K=0.987420882906575
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841082_8.2u  1  2  3  4  PARAMS:
+  Cww=14.15p
+  Rp1=12475
+  Cp1=1.798p
+  Lp1=9.357u
+  Rp2=12475
+  Cp2=1.798p
+  Lp2=9.357u
+  RDC1=0.18
+  RDC2=0.18
+  K=0.988655159492047
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841150_15u  1  2  3  4  PARAMS:
+  Cww=18.34p
+  Rp1=19909
+  Cp1=3.339p
+  Lp1=15.865u
+  Rp2=19909
+  Cp2=3.339p
+  Lp2=15.865u
+  RDC1=0.325
+  RDC2=0.325
+  K=0.990622699787025
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841220_22u  1  2  3  4  PARAMS:
+  Cww=20.85p
+  Rp1=24214
+  Cp1=1.81p
+  Lp1=23.72u
+  Rp2=24214
+  Cp2=1.81p
+  Lp2=23.72u
+  RDC1=0.455
+  RDC2=0.455
+  K=0.990637994609351
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841330_33u  1  2  3  4  PARAMS:
+  Cww=21.63p
+  Rp1=40443
+  Cp1=1.779p
+  Lp1=36.041u
+  Rp2=40443
+  Cp2=1.779p
+  Lp2=36.041u
+  RDC1=0.718
+  RDC2=0.718
+  K=0.990408547473764
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841470_47u  1  2  3  4  PARAMS:
+  Cww=25.4p
+  Rp1=37674
+  Cp1=1.88p
+  Lp1=50.004u
+  Rp2=37674
+  Cp2=1.88p
+  Lp2=50.004u
+  RDC1=0.84
+  RDC2=0.84
+  K=0.990916188997345
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448441100_10u  1  2  3  4  PARAMS:
+  Cww=16.48p
+  Rp1=16318
+  Cp1=1.474p
+  Lp1=13.695u
+  Rp2=16318
+  Cp2=1.474p
+  Lp2=13.695u
+  RDC1=0.21
+  RDC2=0.21
+  K=0.990454441
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_7448841100_10u  1  2  3  4  PARAMS:
+  Cww=16.48p
+  Rp1=16318
+  Cp1=1.474p
+  Lp1=13.695u
+  Rp2=16318
+  Cp2=1.474p
+  Lp2=13.695u
+  RDC1=0.21
+  RDC2=0.21
+  K=0.990454441
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******












