**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMD Power Inductor
* Matchcode:             WE-XHMA
* Library Type:          LTspice
* Version:               rev22b
* Created/modified by:   Ella
* Date and Time:         6/8/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 6030_784393440018_0.18u 1 2
Rp 1 2 393.041
Cp 1 2 5.062p
Rs 1 N3 0.00132
L1 N3 2 0.176u
.ends 6030_784393440018_0.18u
*******
.subckt 6030_784393440033_0.33u 1 2
Rp 1 2 683.781
Cp 1 2 6.324p
Rs 1 N3 0.0021
L1 N3 2 0.316u
.ends 6030_784393440033_0.33u
*******
.subckt 6030_784393440056_0.56u 1 2
Rp 1 2 876.79
Cp 1 2 7.515p
Rs 1 N3 0.0029
L1 N3 2 0.561u
.ends 6030_784393440056_0.56u
*******
.subckt 6030_78439344010_1u 1 2
Rp 1 2 1956
Cp 1 2 7.102p
Rs 1 N3 0.0055
L1 N3 2 1.008u
.ends 6030_78439344010_1u
*******
.subckt 6030_78439344012_1.2u 1 2
Rp 1 2 2178
Cp 1 2 8.182p
Rs 1 N3 0.0064
L1 N3 2 1.105u
.ends 6030_78439344012_1.2u
*******
.subckt 6030_78439344022_2.2u 1 2
Rp 1 2 2927
Cp 1 2 8.36p
Rs 1 N3 0.0105
L1 N3 2 2.182u
.ends 6030_78439344022_2.2u
*******
.subckt 6030_78439344033_3.3u 1 2
Rp 1 2 4970
Cp 1 2 7.979p
Rs 1 N3 0.0192
L1 N3 2 3.247u
.ends 6030_78439344033_3.3u
*******
.subckt 6030_78439344047_4.7u 1 2
Rp 1 2 7211
Cp 1 2 7.002p
Rs 1 N3 0.031
L1 N3 2 4.676u
.ends 6030_78439344047_4.7u
*******
.subckt 6060_78439346047_4.7u 1 2
Rp 1 2 4305
Cp 1 2 7.633p
Rs 1 N3 0.013
L1 N3 2 4.289u
.ends 6060_78439346047_4.7u
*******
.subckt 6060_78439346056_5.6u 1 2
Rp 1 2 5112
Cp 1 2 7.79p
Rs 1 N3 0.015
L1 N3 2 5.311u
.ends 6060_78439346056_5.6u
*******
.subckt 6060_78439346068_6.8u 1 2
Rp 1 2 5867
Cp 1 2 7.976p
Rs 1 N3 0.0176
L1 N3 2 6.553u
.ends 6060_78439346068_6.8u
*******
.subckt 6060_78439346082_8.2u 1 2
Rp 1 2 6820
Cp 1 2 8.668p
Rs 1 N3 0.023
L1 N3 2 7.855u
.ends 6060_78439346082_8.2u
*******
.subckt 6060_78439346100_10u 1 2
Rp 1 2 9786
Cp 1 2 8.192p
Rs 1 N3 0.0265
L1 N3 2 9.539u
.ends 6060_78439346100_10u
*******
.subckt 8080_78439358010_1u 1 2
Rp 1 2 1445
Cp 1 2 8.916p
Rs 1 N3 0.0021
L1 N3 2 1.014u
.ends 8080_78439358010_1u
*******
.subckt 8080_78439358022_2.2u 1 2
Rp 1 2 2282
Cp 1 2 10.434p
Rs 1 N3 0.0037
L1 N3 2 2.209u
.ends 8080_78439358022_2.2u
*******
.subckt 8080_78439358047_4.7u 1 2
Rp 1 2 4439
Cp 1 2 10.924p
Rs 1 N3 0.00865
L1 N3 2 4.785u
.ends 8080_78439358047_4.7u
*******
.subckt 8080_78439358068_6.8u 1 2
Rp 1 2 6545
Cp 1 2 7.924p
Rs 1 N3 0.013
L1 N3 2 6.596u
.ends 8080_78439358068_6.8u
*******
.subckt 8080_78439358100_10u 1 2
Rp 1 2 8417
Cp 1 2 8.116p
Rs 1 N3 0.019
L1 N3 2 10.282u
.ends 8080_78439358100_10u
*******
.subckt 1090_78439369022_2.2u 1 2
Rp 1 2 2074
Cp 1 2 14.601p
Rs 1 N3 0.0022
L1 N3 2 2.242u
.ends 1090_78439369022_2.2u
*******
.subckt 1090_78439369033_3.3u 1 2
Rp 1 2 3017
Cp 1 2 14.697p
Rs 1 N3 0.0034
L1 N3 2 3.164u
.ends 1090_78439369033_3.3u
*******
.subckt 1090_78439369047_4.7u 1 2
Rp 1 2 4114
Cp 1 2 12.704p
Rs 1 N3 0.005
L1 N3 2 4.625u
.ends 1090_78439369047_4.7u
*******
.subckt 1090_78439369056_5.6u 1 2
Rp 1 2 4898
Cp 1 2 13.52p
Rs 1 N3 0.0059
L1 N3 2 5.491u
.ends 1090_78439369056_5.6u
*******
.subckt 1090_78439369068_6.8u 1 2
Rp 1 2 5791
Cp 1 2 14.891p
Rs 1 N3 0.00716
L1 N3 2 7.08u
.ends 1090_78439369068_6.8u
*******
.subckt 1090_78439369082_8.2u 1 2
Rp 1 2 7214
Cp 1 2 12.059p
Rs 1 N3 0.01
L1 N3 2 8.743u
.ends 1090_78439369082_8.2u
*******
.subckt 1090_78439369100_10u 1 2
Rp 1 2 7876
Cp 1 2 13.203p
Rs 1 N3 0.011
L1 N3 2 10.09u
.ends 1090_78439369100_10u
*******
.subckt 1090_78439369150_15u 1 2
Rp 1 2 8204
Cp 1 2 14.622p
Rs 1 N3 0.0148
L1 N3 2 14.546u
.ends 1090_78439369150_15u
*******
.subckt 1510_78439370047_4.7u 1 2
Rp 1 2 4296
Cp 1 2 22.242p
Rs 1 N3 0.0031
L1 N3 2 4.217u
.ends 1510_78439370047_4.7u
*******
.subckt 1510_78439370068_6.8u 1 2
Rp 1 2 5066
Cp 1 2 21.801p
Rs 1 N3 0.0041
L1 N3 2 6.111u
.ends 1510_78439370068_6.8u
*******
.subckt 1510_78439370082_8.2u 1 2
Rp 1 2 6284
Cp 1 2 25.54p
Rs 1 N3 0.0055
L1 N3 2 8.328u
.ends 1510_78439370082_8.2u
*******
.subckt 1510_78439370100_10u 1 2
Rp 1 2 5244
Cp 1 2 29.045p
Rs 1 N3 0.0064
L1 N3 2 10.4u
.ends 1510_78439370100_10u
*******
.subckt 1510_78439370150_15u 1 2
Rp 1 2 7827
Cp 1 2 24.013p
Rs 1 N3 0.0105
L1 N3 2 15.895u
.ends 1510_78439370150_15u
*******
.subckt 1510_78439370220_22u 1 2
Rp 1 2 8204
Cp 1 2 26.195p
Rs 1 N3 0.0125
L1 N3 2 20.695u
.ends 1510_78439370220_22u
*******
.subckt 1510_78439370330_33u 1 2
Rp 1 2 10776
Cp 1 2 27.127p
Rs 1 N3 0.018
L1 N3 2 31.904u
.ends 1510_78439370330_33u
*******
