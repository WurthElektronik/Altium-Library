**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ATG8
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 860010272001_22uF 1 2
Rser 1 3 2.06388553485
Lser 2 4 3.432813032E-09
C1 3 4 0.000022
Rpar 3 4 3333333.33333333
.ends 860010272001_22uF
*******
.subckt 860010272002_33uF 1 2
Rser 1 3 1.64265288281
Lser 2 4 3.113732569E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860010272002_33uF
*******
.subckt 860010272003_47uF 1 2
Rser 1 3 1.30347761752
Lser 2 4 3.668715976E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860010272003_47uF
*******
.subckt 860010272004_68uF 1 2
Rser 1 3 0.879512093366
Lser 2 4 3.972576803E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860010272004_68uF
*******
.subckt 860010272005_100uF 1 2
Rser 1 3 1.03631162149
Lser 2 4 4.359601619E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860010272005_100uF
*******
.subckt 860010272006_120uF 1 2
Rser 1 3 0.857654185063
Lser 2 4 3.643605949E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860010272006_120uF
*******
.subckt 860010272007_150uF 1 2
Rser 1 3 0.610739410975
Lser 2 4 3.980524865E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860010272007_150uF
*******
.subckt 860010273008_180uF 1 2
Rser 1 3 0.41
Lser 2 4 0.00000002
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860010273008_180uF
*******
.subckt 860010273009_220uF 1 2
Rser 1 3 0.399
Lser 2 4 8.576321785E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860010273009_220uF
*******
.subckt 860010273010_330uF 1 2
Rser 1 3 0.26
Lser 2 4 0.0000000203
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860010273010_330uF
*******
.subckt 860010273011_470uF 1 2
Rser 1 3 0.29
Lser 2 4 0.0000000228
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860010273011_470uF
*******
.subckt 860010274012_560uF 1 2
Rser 1 3 0.163
Lser 2 4 0.000000024
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860010274012_560uF
*******
.subckt 860010274013_680uF 1 2
Rser 1 3 0.145
Lser 2 4 0.0000000225
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860010274013_680uF
*******
.subckt 860010274015_1mF 1 2
Rser 1 3 0.205
Lser 2 4 0.0000000232
C1 3 4 0.001
Rpar 3 4 100000
.ends 860010274015_1mF
*******
.subckt 860010275014_820uF 1 2
Rser 1 3 0.122
Lser 2 4 0.0000000252
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860010275014_820uF
*******
.subckt 860010275016_1mF 1 2
Rser 1 3 0.145
Lser 2 4 0.0000000269
C1 3 4 0.001
Rpar 3 4 100000
.ends 860010275016_1mF
*******
.subckt 860010275017_1.2mF 1 2
Rser 1 3 0.092
Lser 2 4 0.0000000225
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860010275017_1.2mF
*******
.subckt 860010275018_1.5mF 1 2
Rser 1 3 0.075
Lser 2 4 0.0000000235
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860010275018_1.5mF
*******
.subckt 860010275019_1.8mF 1 2
Rser 1 3 0.073
Lser 2 4 0.000000025
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860010275019_1.8mF
*******
.subckt 860010275020_2.2mF 1 2
Rser 1 3 0.067
Lser 2 4 0.0000000246
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860010275020_2.2mF
*******
.subckt 860010278021_2.7mF 1 2
Rser 1 3 0.054
Lser 2 4 0.000000024
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860010278021_2.7mF
*******
.subckt 860010278022_3.3mF 1 2
Rser 1 3 0.0504
Lser 2 4 0.0000000268
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860010278022_3.3mF
*******
.subckt 860010278023_3.9mF 1 2
Rser 1 3 0.0335
Lser 2 4 0.000000006
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860010278023_3.9mF
*******
.subckt 860010278024_4.7mF 1 2
Rser 1 3 0.042
Lser 2 4 0.0000000303
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860010278024_4.7mF
*******
.subckt 860010280025_5.6mF 1 2
Rser 1 3 0.041
Lser 2 4 0.0000000334
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860010280025_5.6mF
*******
.subckt 860010280026_6.8mF 1 2
Rser 1 3 0.0385
Lser 2 4 0.0000000329
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860010280026_6.8mF
*******
.subckt 860010280027_8.2mF 1 2
Rser 1 3 0.025
Lser 2 4 0.0000000317
C1 3 4 0.0082
Rpar 3 4 12195.1219512195
.ends 860010280027_8.2mF
*******
.subckt 860010280028_10mF 1 2
Rser 1 3 0.0215
Lser 2 4 0.0000000178
C1 3 4 0.01
Rpar 3 4 10000
.ends 860010280028_10mF
*******
.subckt 860010281029_12mF 1 2
Rser 1 3 0.0175
Lser 2 4 0.0000000086
C1 3 4 0.012
Rpar 3 4 8333.33333333333
.ends 860010281029_12mF
*******
.subckt 860010281030_15mF 1 2
Rser 1 3 0.024
Lser 2 4 0.0000000356
C1 3 4 0.015
Rpar 3 4 6666.66666666667
.ends 860010281030_15mF
*******
.subckt 860010281031_18mF 1 2
Rser 1 3 0.0234
Lser 2 4 0.0000000368
C1 3 4 0.018
Rpar 3 4 5555.55555555556
.ends 860010281031_18mF
*******
.subckt 860010283032_22mF 1 2
Rser 1 3 0.0195
Lser 2 4 0.00000004
C1 3 4 0.022
Rpar 3 4 4545.45454545455
.ends 860010283032_22mF
*******
.subckt 860010283033_33mF 1 2
Rser 1 3 0.0165
Lser 2 4 0.000000035
C1 3 4 0.033
Rpar 3 4 3030.30303030303
.ends 860010283033_33mF
*******
.subckt 860010372001_10uF 1 2
Rser 1 3 2.48763733086
Lser 2 4 4.112727641E-09
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 860010372001_10uF
*******
.subckt 860010372002_22uF 1 2
Rser 1 3 2.27227030586
Lser 2 4 2.874556031E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860010372002_22uF
*******
.subckt 860010372003_33uF 1 2
Rser 1 3 0.78
Lser 2 4 0.0000000085
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860010372003_33uF
*******
.subckt 860010372004_47uF 1 2
Rser 1 3 1.03518743409
Lser 2 4 3.871059877E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860010372004_47uF
*******
.subckt 860010372005_68uF 1 2
Rser 1 3 1.07271061821
Lser 2 4 3.884360416E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860010372005_68uF
*******
.subckt 860010372006_100uF 1 2
Rser 1 3 0.72
Lser 2 4 0.0000000184
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860010372006_100uF
*******
.subckt 860010373007_120uF 1 2
Rser 1 3 0.481131815272
Lser 2 4 4.982100947E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860010373007_120uF
*******
.subckt 860010373008_150uF 1 2
Rser 1 3 0.4002049767
Lser 2 4 4.907053114E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860010373008_150uF
*******
.subckt 860010373009_180uF 1 2
Rser 1 3 0.255
Lser 2 4 0.0000000034
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860010373009_180uF
*******
.subckt 860010373010_220uF 1 2
Rser 1 3 0.29
Lser 2 4 0.0000000238
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860010373010_220uF
*******
.subckt 860010374011_330uF 1 2
Rser 1 3 0.19
Lser 2 4 0.0000000038
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860010374011_330uF
*******
.subckt 860010374012_470uF 1 2
Rser 1 3 0.13
Lser 2 4 0.00000000362
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860010374012_470uF
*******
.subckt 860010374014_680uF 1 2
Rser 1 3 0.135
Lser 2 4 0.0000000312
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860010374014_680uF
*******
.subckt 860010375013_560uF 1 2
Rser 1 3 0.158
Lser 2 4 0.0000000044
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860010375013_560uF
*******
.subckt 860010375015_680uF 1 2
Rser 1 3 0.113
Lser 2 4 0.0000000252
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860010375015_680uF
*******
.subckt 860010375016_820uF 1 2
Rser 1 3 0.103
Lser 2 4 0.0000000244
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860010375016_820uF
*******
.subckt 860010375017_1mF 1 2
Rser 1 3 0.072
Lser 2 4 0.0000000039
C1 3 4 0.001
Rpar 3 4 100000
.ends 860010375017_1mF
*******
.subckt 860010375018_1.2mF 1 2
Rser 1 3 0.081
Lser 2 4 0.0000000288
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860010375018_1.2mF
*******
.subckt 860010375019_1.5mF 1 2
Rser 1 3 0.087
Lser 2 4 0.0000000254
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860010375019_1.5mF
*******
.subckt 860010378020_1.8mF 1 2
Rser 1 3 0.063
Lser 2 4 0.0000000271
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860010378020_1.8mF
*******
.subckt 860010378021_2.2mF 1 2
Rser 1 3 0.04
Lser 2 4 0.000000005
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860010378021_2.2mF
*******
.subckt 860010378022_2.7mF 1 2
Rser 1 3 0.053
Lser 2 4 0.0000000276
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860010378022_2.7mF
*******
.subckt 860010378023_3.3mF 1 2
Rser 1 3 0.038
Lser 2 4 0.00000000596
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860010378023_3.3mF
*******
.subckt 860010380024_3.9mF 1 2
Rser 1 3 0.0419
Lser 2 4 0.0000000297
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860010380024_3.9mF
*******
.subckt 860010380025_4.7mF 1 2
Rser 1 3 0.023
Lser 2 4 0.0000000095
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860010380025_4.7mF
*******
.subckt 860010380026_5.6mF 1 2
Rser 1 3 0.0284
Lser 2 4 0.0000000312
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860010380026_5.6mF
*******
.subckt 860010380027_6.8mF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000337
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860010380027_6.8mF
*******
.subckt 860010380028_8.2mF 1 2
Rser 1 3 0.0265
Lser 2 4 0.000000034
C1 3 4 0.0082
Rpar 3 4 12195.1219512195
.ends 860010380028_8.2mF
*******
.subckt 860010381029_10mF 1 2
Rser 1 3 0.035
Lser 2 4 0.0000000311
C1 3 4 0.01
Rpar 3 4 10000
.ends 860010381029_10mF
*******
.subckt 860010381030_12mF 1 2
Rser 1 3 0.026
Lser 2 4 0.0000000358
C1 3 4 0.012
Rpar 3 4 8333.33333333333
.ends 860010381030_12mF
*******
.subckt 860010383031_15mF 1 2
Rser 1 3 0.02
Lser 2 4 0.000000036
C1 3 4 0.015
Rpar 3 4 6666.66666666667
.ends 860010383031_15mF
*******
.subckt 860010472001_4.7uF 1 2
Rser 1 3 2.50299151711
Lser 2 4 1.736128015E-09
C1 3 4 0.0000047
Rpar 3 4 8333333.33333333
.ends 860010472001_4.7uF
*******
.subckt 860010472002_10uF 1 2
Rser 1 3 1.1
Lser 2 4 0.0000000063
C1 3 4 0.00001
Rpar 3 4 8333333.33333333
.ends 860010472002_10uF
*******
.subckt 860010472003_22uF 1 2
Rser 1 3 1.21755121709
Lser 2 4 4.424663203E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860010472003_22uF
*******
.subckt 860010472004_33uF 1 2
Rser 1 3 1.02973053137
Lser 2 4 4.503431609E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860010472004_33uF
*******
.subckt 860010472005_47uF 1 2
Rser 1 3 1.02887774419
Lser 2 4 3.919583722E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860010472005_47uF
*******
.subckt 860010473006_68uF 1 2
Rser 1 3 0.568501176557
Lser 2 4 4.481745308E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860010473006_68uF
*******
.subckt 860010473007_100uF 1 2
Rser 1 3 0.488708270923
Lser 2 4 4.372078024E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860010473007_100uF
*******
.subckt 860010473008_120uF 1 2
Rser 1 3 0.308
Lser 2 4 0.0000000029
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860010473008_120uF
*******
.subckt 860010473009_150uF 1 2
Rser 1 3 0.275
Lser 2 4 0.0000000188
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860010473009_150uF
*******
.subckt 860010473010_180uF 1 2
Rser 1 3 0.26
Lser 2 4 0.0000000028
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860010473010_180uF
*******
.subckt 860010473011_220uF 1 2
Rser 1 3 0.2
Lser 2 4 0.0000000024
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860010473011_220uF
*******
.subckt 860010474012_330uF 1 2
Rser 1 3 0.15
Lser 2 4 0.0000000036
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860010474012_330uF
*******
.subckt 860010474013_470uF 1 2
Rser 1 3 0.118
Lser 2 4 0.000000003
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860010474013_470uF
*******
.subckt 860010475014_560uF 1 2
Rser 1 3 0.118
Lser 2 4 0.000000004
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860010475014_560uF
*******
.subckt 860010475015_680uF 1 2
Rser 1 3 0.093
Lser 2 4 0.000000004
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860010475015_680uF
*******
.subckt 860010475016_820uF 1 2
Rser 1 3 0.088
Lser 2 4 0.0000000237
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860010475016_820uF
*******
.subckt 860010475017_1mF 1 2
Rser 1 3 0.063
Lser 2 4 0.0000000255
C1 3 4 0.001
Rpar 3 4 100000
.ends 860010475017_1mF
*******
.subckt 860010478018_1.2mF 1 2
Rser 1 3 0.086
Lser 2 4 0.0000000278
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860010478018_1.2mF
*******
.subckt 860010478019_1.5mF 1 2
Rser 1 3 0.073
Lser 2 4 0.0000000268
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860010478019_1.5mF
*******
.subckt 860010478020_1.8mF 1 2
Rser 1 3 0.055
Lser 2 4 0.0000000258
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860010478020_1.8mF
*******
.subckt 860010478021_2.2mF 1 2
Rser 1 3 0.048
Lser 2 4 0.000000029
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860010478021_2.2mF
*******
.subckt 860010480022_2.7mF 1 2
Rser 1 3 0.035
Lser 2 4 0.0000000298
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860010480022_2.7mF
*******
.subckt 860010480023_3.3mF 1 2
Rser 1 3 0.035
Lser 2 4 0.000000029
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860010480023_3.3mF
*******
.subckt 860010480024_3.9mF 1 2
Rser 1 3 0.028
Lser 2 4 0.0000000328
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860010480024_3.9mF
*******
.subckt 860010480025_4.7mF 1 2
Rser 1 3 0.029
Lser 2 4 0.0000000375
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860010480025_4.7mF
*******
.subckt 860010481026_5.6mF 1 2
Rser 1 3 0.027
Lser 2 4 0.0000000323
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860010481026_5.6mF
*******
.subckt 860010481027_6.8mF 1 2
Rser 1 3 0.0255
Lser 2 4 0.0000000348
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860010481027_6.8mF
*******
.subckt 860010481028_8.2mF 1 2
Rser 1 3 0.024
Lser 2 4 0.0000000306
C1 3 4 0.0082
Rpar 3 4 12195.1219512195
.ends 860010481028_8.2mF
*******
.subckt 860010483029_10mF 1 2
Rser 1 3 0.0225
Lser 2 4 0.0000000412
C1 3 4 0.01
Rpar 3 4 10000
.ends 860010483029_10mF
*******
.subckt 860010572001_4.7uF 1 2
Rser 1 3 1.17
Lser 2 4 0.000000007
C1 3 4 0.0000047
Rpar 3 4 11666666.6666667
.ends 860010572001_4.7uF
*******
.subckt 860010572002_10uF 1 2
Rser 1 3 2.6734604472
Lser 2 4 1.683206479E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860010572002_10uF
*******
.subckt 860010572003_22uF 1 2
Rser 1 3 0.97915012213
Lser 2 4 4.327727353E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 860010572003_22uF
*******
.subckt 860010572004_33uF 1 2
Rser 1 3 0.81881047648
Lser 2 4 4.592522954E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860010572004_33uF
*******
.subckt 860010572005_47uF 1 2
Rser 1 3 0.896216410917
Lser 2 4 0.000000003276938
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860010572005_47uF
*******
.subckt 860010573006_68uF 1 2
Rser 1 3 0.456922433265
Lser 2 4 4.281681279E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860010573006_68uF
*******
.subckt 860010573007_100uF 1 2
Rser 1 3 0.38
Lser 2 4 0.00000000298
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860010573007_100uF
*******
.subckt 860010574008_120uF 1 2
Rser 1 3 0.40147327634
Lser 2 4 4.642502404E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860010574008_120uF
*******
.subckt 860010574009_150uF 1 2
Rser 1 3 0.4
Lser 2 4 0.0000000145
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860010574009_150uF
*******
.subckt 860010574010_180uF 1 2
Rser 1 3 0.225
Lser 2 4 0.0000000034
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860010574010_180uF
*******
.subckt 860010574011_220uF 1 2
Rser 1 3 0.19
Lser 2 4 0.0000000037
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860010574011_220uF
*******
.subckt 860010575012_330uF 1 2
Rser 1 3 0.185
Lser 2 4 0.0000000308
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860010575012_330uF
*******
.subckt 860010575013_470uF 1 2
Rser 1 3 0.073
Lser 2 4 0.00000000396
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860010575013_470uF
*******
.subckt 860010575014_560uF 1 2
Rser 1 3 0.087
Lser 2 4 0.0000000276
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860010575014_560uF
*******
.subckt 860010575015_680uF 1 2
Rser 1 3 0.082
Lser 2 4 0.0000000275
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860010575015_680uF
*******
.subckt 860010578016_820uF 1 2
Rser 1 3 0.081
Lser 2 4 0.0000000259
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860010578016_820uF
*******
.subckt 860010578017_1mF 1 2
Rser 1 3 0.064
Lser 2 4 0.0000000055
C1 3 4 0.001
Rpar 3 4 100000
.ends 860010578017_1mF
*******
.subckt 860010578018_1.2mF 1 2
Rser 1 3 0.062
Lser 2 4 0.0000000055
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860010578018_1.2mF
*******
.subckt 860010578019_1.5mF 1 2
Rser 1 3 0.0505
Lser 2 4 0.0000000299
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860010578019_1.5mF
*******
.subckt 860010580020_1.8mF 1 2
Rser 1 3 0.039
Lser 2 4 0.0000000289
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860010580020_1.8mF
*******
.subckt 860010580021_2.2mF 1 2
Rser 1 3 0.0265
Lser 2 4 0.0000000096
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860010580021_2.2mF
*******
.subckt 860010580022_2.7mF 1 2
Rser 1 3 0.023
Lser 2 4 0.0000000078
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860010580022_2.7mF
*******
.subckt 860010580023_3.3mF 1 2
Rser 1 3 0.0275
Lser 2 4 0.0000000102
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860010580023_3.3mF
*******
.subckt 860010581024_3.9mF 1 2
Rser 1 3 0.025
Lser 2 4 0.00000000796
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860010581024_3.9mF
*******
.subckt 860010581025_4.7mF 1 2
Rser 1 3 0.026
Lser 2 4 0.000000031
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860010581025_4.7mF
*******
.subckt 860010581026_5.6mF 1 2
Rser 1 3 0.026
Lser 2 4 0.0000000338
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860010581026_5.6mF
*******
.subckt 860010583027_6.8mF 1 2
Rser 1 3 0.022
Lser 2 4 0.0000000352
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860010583027_6.8mF
*******
.subckt 860010672001_100nF 1 2
Rser 1 3 3.09403328355
Lser 2 4 3.756071489E-09
C1 3 4 0.0000001
Rpar 3 4 16666666.6666667
.ends 860010672001_100nF
*******
.subckt 860010672002_220nF 1 2
Rser 1 3 2.7030039461
Lser 2 4 2.814543386E-09
C1 3 4 0.00000022
Rpar 3 4 16666666.6666667
.ends 860010672002_220nF
*******
.subckt 860010672003_330nF 1 2
Rser 1 3 1.55
Lser 2 4 1.31745210618708E-07
C1 3 4 0.00000033
Rpar 3 4 16666666.6666667
.ends 860010672003_330nF
*******
.subckt 860010672004_470nF 1 2
Rser 1 3 2.6630641601
Lser 2 4 3.418092208E-09
C1 3 4 0.00000047
Rpar 3 4 16666666.6666667
.ends 860010672004_470nF
*******
.subckt 860010672005_1uF 1 2
Rser 1 3 3.02266243136
Lser 2 4 4.262975117E-09
C1 3 4 0.000001
Rpar 3 4 16666666.6666667
.ends 860010672005_1uF
*******
.subckt 860010672006_2.2uF 1 2
Rser 1 3 2.44273654792
Lser 2 4 1.706914429E-09
C1 3 4 0.0000022
Rpar 3 4 16666666.6666667
.ends 860010672006_2.2uF
*******
.subckt 860010672007_3.3uF 1 2
Rser 1 3 0.86
Lser 2 4 0.0000000059
C1 3 4 0.0000033
Rpar 3 4 16666666.6666667
.ends 860010672007_3.3uF
*******
.subckt 860010672008_4.7uF 1 2
Rser 1 3 2.4290928933
Lser 2 4 4.037180944E-09
C1 3 4 0.0000047
Rpar 3 4 16666666.6666667
.ends 860010672008_4.7uF
*******
.subckt 860010672009_10uF 1 2
Rser 1 3 1.91533261427
Lser 2 4 3.377044238E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860010672009_10uF
*******
.subckt 860010672010_22uF 1 2
Rser 1 3 0.785920274015
Lser 2 4 5.463190311E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860010672010_22uF
*******
.subckt 860010672011_33uF 1 2
Rser 1 3 0.51
Lser 2 4 0.0000000057
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860010672011_33uF
*******
.subckt 860010673012_47uF 1 2
Rser 1 3 0.625207993849
Lser 2 4 4.314152653E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860010673012_47uF
*******
.subckt 860010674013_68uF 1 2
Rser 1 3 0.275
Lser 2 4 0.0000000075
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860010674013_68uF
*******
.subckt 860010674014_100uF 1 2
Rser 1 3 0.278
Lser 2 4 0.0000000033
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860010674014_100uF
*******
.subckt 860010674015_120uF 1 2
Rser 1 3 0.245
Lser 2 4 0.0000000244
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860010674015_120uF
*******
.subckt 860010675016_150uF 1 2
Rser 1 3 0.32
Lser 2 4 0.0000000225
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860010675016_150uF
*******
.subckt 860010675017_180uF 1 2
Rser 1 3 0.353780164787
Lser 2 4 5.088657592E-09
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860010675017_180uF
*******
.subckt 860010675018_220uF 1 2
Rser 1 3 0.255
Lser 2 4 0.0000000218
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860010675018_220uF
*******
.subckt 860010675019_330uF 1 2
Rser 1 3 0.137
Lser 2 4 0.0000000203
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860010675019_330uF
*******
.subckt 860010675020_470uF 1 2
Rser 1 3 0.085
Lser 2 4 0.0000000034
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860010675020_470uF
*******
.subckt 860010678021_560uF 1 2
Rser 1 3 0.0805
Lser 2 4 0.0000000262
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860010678021_560uF
*******
.subckt 860010678022_680uF 1 2
Rser 1 3 0.064
Lser 2 4 0.0000000056
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860010678022_680uF
*******
.subckt 860010678023_820uF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000063
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860010678023_820uF
*******
.subckt 860010678024_1mF 1 2
Rser 1 3 0.057
Lser 2 4 0.0000000272
C1 3 4 0.001
Rpar 3 4 100000
.ends 860010678024_1mF
*******
.subckt 860010680025_1.2mF 1 2
Rser 1 3 0.069
Lser 2 4 0.0000000291
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860010680025_1.2mF
*******
.subckt 860010680026_1.5mF 1 2
Rser 1 3 0.054
Lser 2 4 0.0000000315
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860010680026_1.5mF
*******
.subckt 860010680027_1.8mF 1 2
Rser 1 3 0.0515
Lser 2 4 0.0000000288
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860010680027_1.8mF
*******
.subckt 860010680028_2.2mF 1 2
Rser 1 3 0.026
Lser 2 4 0.0000000076
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860010680028_2.2mF
*******
.subckt 860010681029_2.7mF 1 2
Rser 1 3 0.0495
Lser 2 4 0.0000000348
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860010681029_2.7mF
*******
.subckt 860010681030_3.3mF 1 2
Rser 1 3 0.0285
Lser 2 4 0.0000000364
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860010681030_3.3mF
*******
.subckt 860010681031_3.9mF 1 2
Rser 1 3 0.0366
Lser 2 4 0.0000000338
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860010681031_3.9mF
*******
.subckt 860010683032_4.7mF 1 2
Rser 1 3 0.015
Lser 2 4 0.0000000097
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860010683032_4.7mF
*******
.subckt 860010772001_100nF 1 2
Rser 1 3 2.89490999071
Lser 2 4 3.019562708E-09
C1 3 4 0.0000001
Rpar 3 4 21000000
.ends 860010772001_100nF
*******
.subckt 860010772002_220nF 1 2
Rser 1 3 2.72154827867
Lser 2 4 2.899519755E-09
C1 3 4 0.00000022
Rpar 3 4 21000000
.ends 860010772002_220nF
*******
.subckt 860010772003_330nF 1 2
Rser 1 3 1.90260444906
Lser 2 4 3.267853108E-09
C1 3 4 0.00000033
Rpar 3 4 21000000
.ends 860010772003_330nF
*******
.subckt 860010772004_470nF 1 2
Rser 1 3 2.59135105628
Lser 2 4 3.170337084E-09
C1 3 4 0.00000047
Rpar 3 4 21000000
.ends 860010772004_470nF
*******
.subckt 860010772005_1uF 1 2
Rser 1 3 1.9
Lser 2 4 5.874602569E-09
C1 3 4 0.000001
Rpar 3 4 21000000
.ends 860010772005_1uF
*******
.subckt 860010772006_2.2uF 1 2
Rser 1 3 0.95
Lser 2 4 0.000000007
C1 3 4 0.0000022
Rpar 3 4 21000000
.ends 860010772006_2.2uF
*******
.subckt 860010772007_3.3uF 1 2
Rser 1 3 2.2052715946
Lser 2 4 3.191475815E-09
C1 3 4 0.0000033
Rpar 3 4 21000000
.ends 860010772007_3.3uF
*******
.subckt 860010772008_4.7uF 1 2
Rser 1 3 1.39380961103
Lser 2 4 3.361147757E-09
C1 3 4 0.0000047
Rpar 3 4 21000000
.ends 860010772008_4.7uF
*******
.subckt 860010772009_10uF 1 2
Rser 1 3 1.05
Lser 2 4 0.0000000061
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860010772009_10uF
*******
.subckt 860010773010_22uF 1 2
Rser 1 3 1.51868187584
Lser 2 4 3.418279081E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860010773010_22uF
*******
.subckt 860010773011_33uF 1 2
Rser 1 3 1.0006070562
Lser 2 4 3.985238411E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860010773011_33uF
*******
.subckt 860010773012_47uF 1 2
Rser 1 3 0.55978172043
Lser 2 4 3.875005269E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860010773012_47uF
*******
.subckt 860010774013_68uF 1 2
Rser 1 3 0.21
Lser 2 4 0.000000008
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860010774013_68uF
*******
.subckt 860010775014_100uF 1 2
Rser 1 3 0.33
Lser 2 4 0.00000000386
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860010775014_100uF
*******
.subckt 860010775015_120uF 1 2
Rser 1 3 0.149
Lser 2 4 0.0000000216
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860010775015_120uF
*******
.subckt 860010775016_150uF 1 2
Rser 1 3 0.129
Lser 2 4 0.0000000246
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860010775016_150uF
*******
.subckt 860010775017_180uF 1 2
Rser 1 3 0.077
Lser 2 4 0.00000000455
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860010775017_180uF
*******
.subckt 860010775018_220uF 1 2
Rser 1 3 0.067
Lser 2 4 0.0000000041
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860010775018_220uF
*******
.subckt 860010775019_330uF 1 2
Rser 1 3 0.135
Lser 2 4 0.0000000138
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860010775019_330uF
*******
.subckt 860010778020_470uF 1 2
Rser 1 3 0.072
Lser 2 4 0.0000000245
C1 3 4 0.00047
Rpar 3 4 212765.957446808
.ends 860010778020_470uF
*******
.subckt 860010778021_560uF 1 2
Rser 1 3 0.06
Lser 2 4 0.0000000301
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860010778021_560uF
*******
.subckt 860010780022_680uF 1 2
Rser 1 3 0.04
Lser 2 4 0.000000031
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860010780022_680uF
*******
.subckt 860010780023_820uF 1 2
Rser 1 3 0.04
Lser 2 4 0.0000000308
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860010780023_820uF
*******
.subckt 860010780024_1mF 1 2
Rser 1 3 0.041
Lser 2 4 0.0000000299
C1 3 4 0.001
Rpar 3 4 100000
.ends 860010780024_1mF
*******
.subckt 860010780025_1.2mF 1 2
Rser 1 3 0.034
Lser 2 4 0.0000000354
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860010780025_1.2mF
*******
.subckt 860010780026_1.5mF 1 2
Rser 1 3 0.032
Lser 2 4 0.0000000319
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860010780026_1.5mF
*******
.subckt 860010780027_1.8mF 1 2
Rser 1 3 0.0278
Lser 2 4 0.0000000325
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860010780027_1.8mF
*******
.subckt 860010781028_2.2mF 1 2
Rser 1 3 0.0195
Lser 2 4 0.0000000083
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860010781028_2.2mF
*******
.subckt 860010783029_2.7mF 1 2
Rser 1 3 0.023
Lser 2 4 0.000000034
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860010783029_2.7mF
*******
.subckt 860010783030_3.3mF 1 2
Rser 1 3 0.024
Lser 2 4 2.2553928962E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860010783030_3.3mF
*******
.subckt 860011373001_470nF 1 2
Rser 1 3 1.58338764937
Lser 2 4 4.691742076E-09
C1 3 4 0.00000047
Rpar 3 4 133333333.333333
.ends 860011373001_470nF
*******
.subckt 860011373002_1uF 1 2
Rser 1 3 1.3713972414
Lser 2 4 3.538082107E-09
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 860011373002_1uF
*******
.subckt 860011374003_2.2uF 1 2
Rser 1 3 1.32124878641
Lser 2 4 4.291371163E-09
C1 3 4 0.0000022
Rpar 3 4 45454545.4545455
.ends 860011374003_2.2uF
*******
.subckt 860011374004_3.3uF 1 2
Rser 1 3 1.0892554435
Lser 2 4 3.781643523E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 860011374004_3.3uF
*******
.subckt 860011374005_4.7uF 1 2
Rser 1 3 1.07032089826
Lser 2 4 5.304520543E-09
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 860011374005_4.7uF
*******
.subckt 860011375006_10uF 1 2
Rser 1 3 0.69785201933
Lser 2 4 4.233915002E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860011375006_10uF
*******
.subckt 860011378007_22uF 1 2
Rser 1 3 0.674269667594
Lser 2 4 6.680332811E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860011378007_22uF
*******
.subckt 860011378008_33uF 1 2
Rser 1 3 0.595
Lser 2 4 1.0849880001E-08
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860011378008_33uF
*******
.subckt 860011380009_47uF 1 2
Rser 1 3 0.567572175543
Lser 2 4 1.1756797098E-08
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860011380009_47uF
*******
.subckt 860011380010_68uF 1 2
Rser 1 3 0.496289860705
Lser 2 4 1.1249087065E-08
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860011380010_68uF
*******
.subckt 860011381011_68uF 1 2
Rser 1 3 0.510234849282
Lser 2 4 1.2049123149E-08
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860011381011_68uF
*******
.subckt 860011381012_100uF 1 2
Rser 1 3 0.406664090715
Lser 2 4 1.2913173134E-08
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860011381012_100uF
*******
.subckt 860011381013_120uF 1 2
Rser 1 3 0.422719278176
Lser 2 4 1.1401288119E-08
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860011381013_120uF
*******
