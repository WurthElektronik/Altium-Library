**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Wire Wound Inductor 
* Matchcode:              WE-GF 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-08
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1210_744764002_0.22u 1 2
Rp 1 2 1601.45
Cp 1 2 0.236p
Rs 1 N3 0.32
L1 N3 2 0.22u
.ends 1210_744764002_0.22u
*******
.subckt 1210_7447640027_0.27u 1 2
Rp 1 2 1923.55
Cp 1 2 0.253p
Rs 1 N3 0.36
L1 N3 2 0.27u
.ends 1210_7447640027_0.27u
*******
.subckt 1210_744764003_0.39u 1 2
Rp 1 2 2681.26
Cp 1 2 0.231p
Rs 1 N3 0.45
L1 N3 2 0.39u
.ends 1210_744764003_0.39u
*******
.subckt 1210_7447640033_0.33u 1 2
Rp 1 2 2267.35
Cp 1 2 0.239p
Rs 1 N3 0.4
L1 N3 2 0.33u
.ends 1210_7447640033_0.33u
*******
.subckt 1210_744764004_0.47u 1 2
Rp 1 2 3340.08
Cp 1 2 0.219p
Rs 1 N3 0.5
L1 N3 2 0.47u
.ends 1210_744764004_0.47u
*******
.subckt 1210_744764005_0.56u 1 2
Rp 1 2 4322.04
Cp 1 2 0.216p
Rs 1 N3 0.55
L1 N3 2 0.56u
.ends 1210_744764005_0.56u
*******
.subckt 1210_744764006_0.68u 1 2
Rp 1 2 5213.16
Cp 1 2 0.214p
Rs 1 N3 0.6
L1 N3 2 0.68u
.ends 1210_744764006_0.68u
*******
.subckt 1210_7447640082_0.82u 1 2
Rp 1 2 5392.96
Cp 1 2 0.197p
Rs 1 N3 0.65
L1 N3 2 0.82u
.ends 1210_7447640082_0.82u
*******
.subckt 1210_74476401_1u 1 2
Rp 1 2 4264.75
Cp 1 2 0.196p
Rs 1 N3 0.7
L1 N3 2 1u
.ends 1210_74476401_1u
*******
.subckt 1210_744764012_1.2u 1 2
Rp 1 2 5359.84
Cp 1 2 0.223p
Rs 1 N3 0.75
L1 N3 2 1.2u
.ends 1210_744764012_1.2u
*******
.subckt 1210_744764015_1.5u 1 2
Rp 1 2 5198.78
Cp 1 2 0.291p
Rs 1 N3 0.85
L1 N3 2 1.5u
.ends 1210_744764015_1.5u
*******
.subckt 1210_744764018_1.8u 1 2
Rp 1 2 6371.37
Cp 1 2 0.433p
Rs 1 N3 0.9
L1 N3 2 1.8u
.ends 1210_744764018_1.8u
*******
.subckt 1210_74476402_2.2u 1 2
Rp 1 2 7534.54
Cp 1 2 0.66p
Rs 1 N3 1
L1 N3 2 2.2u
.ends 1210_74476402_2.2u
*******
.subckt 1210_744764027_2.7u 1 2
Rp 1 2 7615.94
Cp 1 2 1.007p
Rs 1 N3 1.1
L1 N3 2 2.7u
.ends 1210_744764027_2.7u
*******
.subckt 1210_74476403_3.3u 1 2
Rp 1 2 8923.53
Cp 1 2 1.456p
Rs 1 N3 1.2
L1 N3 2 3.3u
.ends 1210_74476403_3.3u
*******
.subckt 1210_744764039_3.9u 1 2
Rp 1 2 10290.6
Cp 1 2 1.635p
Rs 1 N3 1.3
L1 N3 2 3.9u
.ends 1210_744764039_3.9u
*******
.subckt 1210_74476404_4.7u 1 2
Rp 1 2 12188.3
Cp 1 2 1.664p
Rs 1 N3 1.5
L1 N3 2 4.7u
.ends 1210_74476404_4.7u
*******
.subckt 1210_74476406_6.8u 1 2
Rp 1 2 16570.2
Cp 1 2 1.677p
Rs 1 N3 1.8
L1 N3 2 6.8u
.ends 1210_74476406_6.8u
*******
.subckt 1210_74476410_10u 1 2
Rp 1 2 27227.9
Cp 1 2 1.532p
Rs 1 N3 2.1
L1 N3 2 10u
.ends 1210_74476410_10u
*******
.subckt 1210_744764112_12u 1 2
Rp 1 2 29691.4
Cp 1 2 1.623p
Rs 1 N3 2.5
L1 N3 2 12u
.ends 1210_744764112_12u
*******
.subckt 1210_744764115_15u 1 2
Rp 1 2 37035.7
Cp 1 2 1.824p
Rs 1 N3 2.8
L1 N3 2 15u
.ends 1210_744764115_15u
*******
.subckt 1210_744764118_18u 1 2
Rp 1 2 57729.2
Cp 1 2 1.668p
Rs 1 N3 3.3
L1 N3 2 18u
.ends 1210_744764118_18u
*******
.subckt 1210_744764122_22u 1 2
Rp 1 2 97573.1
Cp 1 2 1.768p
Rs 1 N3 3.7
L1 N3 2 22u
.ends 1210_744764122_22u
*******
.subckt 1210_744764133_33u 1 2
Rp 1 2 391578
Cp 1 2 1.8p
Rs 1 N3 5.6
L1 N3 2 33u
.ends 1210_744764133_33u
*******
.subckt 1210_744764139_39u 1 2
Rp 1 2 495039
Cp 1 2 1.758p
Rs 1 N3 6.4
L1 N3 2 39u
.ends 1210_744764139_39u
*******
.subckt 1210_744764147_47u 1 2
Rp 1 2 462536
Cp 1 2 1.83p
Rs 1 N3 7
L1 N3 2 47u
.ends 1210_744764147_47u
*******
.subckt 1210_744764156_56u 1 2
Rp 1 2 349813
Cp 1 2 1.713p
Rs 1 N3 8
L1 N3 2 56u
.ends 1210_744764156_56u
*******
.subckt 1210_744764168_68u 1 2
Rp 1 2 277653
Cp 1 2 1.862p
Rs 1 N3 9
L1 N3 2 68u
.ends 1210_744764168_68u
*******
.subckt 1210_74476420_100u 1 2
Rp 1 2 2110000
Cp 1 2 1.754p
Rs 1 N3 11
L1 N3 2 100u
.ends 1210_74476420_100u
*******
.subckt 1812_744766001_0.1u 1 2
Rp 1 2 781.599
Cp 1 2 0.365p
Rs 1 N3 0.44
L1 N3 2 0.1u
.ends 1812_744766001_0.1u
*******
.subckt 1812_7447660033_0.33u 1 2
Rp 1 2 2481.32
Cp 1 2 0.324p
Rs 1 N3 0.4
L1 N3 2 0.33u
.ends 1812_7447660033_0.33u
*******
.subckt 1812_7447660039_0.39u 1 2
Rp 1 2 1449.41
Cp 1 2 0.719p
Rs 1 N3 0.45
L1 N3 2 0.39u
.ends 1812_7447660039_0.39u
*******
.subckt 1812_7447660068_0.68u 1 2
Rp 1 2 4624.6
Cp 1 2 0.359p
Rs 1 N3 0.6
L1 N3 2 0.68u
.ends 1812_7447660068_0.68u
*******
.subckt 1812_7447660082_0.82u 1 2
Rp 1 2 5111.41
Cp 1 2 0.353p
Rs 1 N3 0.67
L1 N3 2 0.82u
.ends 1812_7447660082_0.82u
*******
.subckt 1812_74476601_1u 1 2
Rp 1 2 3733.08
Cp 1 2 0.327p
Rs 1 N3 0.5
L1 N3 2 1u
.ends 1812_74476601_1u
*******
.subckt 1812_744766012_1.2u 1 2
Rp 1 2 4330.43
Cp 1 2 0.323p
Rs 1 N3 0.55
L1 N3 2 1.2u
.ends 1812_744766012_1.2u
*******
.subckt 1812_744766015_1.5u 1 2
Rp 1 2 5144.67
Cp 1 2 0.308p
Rs 1 N3 0.6
L1 N3 2 1.5u
.ends 1812_744766015_1.5u
*******
.subckt 1812_744766018_1.8u 1 2
Rp 1 2 6426.75
Cp 1 2 0.301p
Rs 1 N3 0.65
L1 N3 2 1.8u
.ends 1812_744766018_1.8u
*******
.subckt 1812_74476602_2.2u 1 2
Rp 1 2 7094.39
Cp 1 2 0.304p
Rs 1 N3 0.7
L1 N3 2 2.2u
.ends 1812_74476602_2.2u
*******
.subckt 1812_74476603_3.3u 1 2
Rp 1 2 11019.3
Cp 1 2 0.463p
Rs 1 N3 0.8
L1 N3 2 3.3u
.ends 1812_74476603_3.3u
*******
.subckt 1812_744766039_3.9u 1 2
Rp 1 2 10686.4
Cp 1 2 0.75p
Rs 1 N3 0.9
L1 N3 2 3.9u
.ends 1812_744766039_3.9u
*******
.subckt 1812_74476604_4.7u 1 2
Rp 1 2 13001.6
Cp 1 2 1.007p
Rs 1 N3 1
L1 N3 2 4.7u
.ends 1812_74476604_4.7u
*******
.subckt 1812_744766056_5.6u 1 2
Rp 1 2 12846.1
Cp 1 2 1.213p
Rs 1 N3 1.1
L1 N3 2 5.6u
.ends 1812_744766056_5.6u
*******
.subckt 1812_74476606_6.8u 1 2
Rp 1 2 13128.4
Cp 1 2 1.816p
Rs 1 N3 1.2
L1 N3 2 6.8u
.ends 1812_74476606_6.8u
*******
.subckt 1812_744766082_8.2u 1 2
Rp 1 2 8556.2
Cp 1 2 5.351p
Rs 1 N3 1.4
L1 N3 2 8.2u
.ends 1812_744766082_8.2u
*******
.subckt 1812_74476610_10u 1 2
Rp 1 2 29635.4
Cp 1 2 3.281p
Rs 1 N3 1.6
L1 N3 2 10u
.ends 1812_74476610_10u
*******
.subckt 1812_744766115_15u 1 2
Rp 1 2 39780.5
Cp 1 2 2.671p
Rs 1 N3 2.5
L1 N3 2 15u
.ends 1812_744766115_15u
*******
.subckt 1812_744766118_18u 1 2
Rp 1 2 45623.8
Cp 1 2 3.252p
Rs 1 N3 2.8
L1 N3 2 18u
.ends 1812_744766118_18u
*******
.subckt 1812_744766122_22u 1 2
Rp 1 2 61782.9
Cp 1 2 2.867p
Rs 1 N3 3.2
L1 N3 2 22u
.ends 1812_744766122_22u
*******
.subckt 1812_744766133_33u 1 2
Rp 1 2 101942
Cp 1 2 3.179p
Rs 1 N3 4
L1 N3 2 33u
.ends 1812_744766133_33u
*******
.subckt 1812_744766147_47u 1 2
Rp 1 2 161500
Cp 1 2 3.693p
Rs 1 N3 5
L1 N3 2 47u
.ends 1812_744766147_47u
*******
.subckt 1812_744766156_56u 1 2
Rp 1 2 51733.6
Cp 1 2 6.494p
Rs 1 N3 5.5
L1 N3 2 56u
.ends 1812_744766156_56u
*******
.subckt 1812_744766168_68u 1 2
Rp 1 2 59107.8
Cp 1 2 6.747p
Rs 1 N3 6
L1 N3 2 68u
.ends 1812_744766168_68u
*******
.subckt 1812_74476620_100u 1 2
Rp 1 2 5074.4
Cp 1 2 3.101p
Rs 1 N3 8
L1 N3 2 100u
.ends 1812_74476620_100u
*******
.subckt 1812_744766215_150u 1 2
Rp 1 2 177652
Cp 1 2 2.818p
Rs 1 N3 9
L1 N3 2 150u
.ends 1812_744766215_150u
*******
.subckt 1812_744766218_180u 1 2
Rp 1 2 437287
Cp 1 2 2.532p
Rs 1 N3 9.5
L1 N3 2 180u
.ends 1812_744766218_180u
*******
.subckt 1812_744766220_220u 1 2
Rp 1 2 404577
Cp 1 2 2.481p
Rs 1 N3 10
L1 N3 2 220u
.ends 1812_744766220_220u
*******
.subckt 1812_744766233_330u 1 2
Rp 1 2 664486
Cp 1 2 2.594p
Rs 1 N3 14
L1 N3 2 330u
.ends 1812_744766233_330u
*******
.subckt 1812_744766239_390u 1 2
Rp 1 2 377818
Cp 1 2 2.571p
Rs 1 N3 18
L1 N3 2 390u
.ends 1812_744766239_390u
*******
.subckt 1812_74476624_470u 1 2
Rp 1 2 165751
Cp 1 2 5.389p
Rs 1 N3 26
L1 N3 2 470u
.ends 1812_74476624_470u
*******
.subckt 1812_74476625_560u 1 2
Rp 1 2 179770
Cp 1 2 5.795p
Rs 1 N3 30
L1 N3 2 560u
.ends 1812_74476625_560u
*******
.subckt 1812_74476626_680u 1 2
Rp 1 2 368030
Cp 1 2 2.953p
Rs 1 N3 30
L1 N3 2 680u
.ends 1812_74476626_680u
*******
.subckt 1812_74476628_820u 1 2
Rp 1 2 230154
Cp 1 2 5.036p
Rs 1 N3 45
L1 N3 2 820u
.ends 1812_74476628_820u
*******
.subckt 1812_74476630_1m 1 2
Rp 1 2 112994
Cp 1 2 2.739p
Rs 1 N3 50
L1 N3 2 1000u
.ends 1812_74476630_1m
*******
