**************************************************
* Manufacturer:          Würth Elektronik
* Kinds:                 Shielded Power Inductor
* Matchcode:             WE-XHMI
* Library Type:          LTspice
* Version:               rev24a
* Created/modified by:   Ella
* Date and Time:         01/10/2024
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2024 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1090_74439369015_1.5u 1 2
Rp 1 2 1195
Cp 1 2 19.206p
Rs 1 N3 0.00146
L1 N3 2 1.349u
.ends 1090_74439369015_1.5u
*******
.subckt 1090_74439369022_2.2u 1 2
Rp 1 2 2074
Cp 1 2 14.601p
Rs 1 N3 0.0022
L1 N3 2 2.242u
.ends 1090_74439369022_2.2u
*******
.subckt 1090_74439369033_3.3u 1 2
Rp 1 2 3017
Cp 1 2 14.697p
Rs 1 N3 0.0034
L1 N3 2 3.164u
.ends 1090_74439369033_3.3u
*******
.subckt 1090_74439369047_4.7u 1 2
Rp 1 2 4114
Cp 1 2 12.704p
Rs 1 N3 0.005
L1 N3 2 4.625u
.ends 1090_74439369047_4.7u
*******
.subckt 1090_74439369056_5.6u 1 2
Rp 1 2 4898
Cp 1 2 13.52p
Rs 1 N3 0.0059
L1 N3 2 5.491u
.ends 1090_74439369056_5.6u
*******
.subckt 1090_74439369068_6.8u 1 2
Rp 1 2 5791
Cp 1 2 14.891p
Rs 1 N3 0.00716
L1 N3 2 7.08u
.ends 1090_74439369068_6.8u
*******
.subckt 1090_74439369082_8.2u 1 2
Rp 1 2 7214
Cp 1 2 12.059p
Rs 1 N3 0.01
L1 N3 2 8.743u
.ends 1090_74439369082_8.2u
*******
.subckt 1090_74439369100_10u 1 2
Rp 1 2 7876
Cp 1 2 13.203p
Rs 1 N3 0.011
L1 N3 2 10.09u
.ends 1090_74439369100_10u
*******
.subckt 1090_74439369150_15u 1 2
Rp 1 2 8204
Cp 1 2 14.622p
Rs 1 N3 0.0148
L1 N3 2 14.546u
.ends 1090_74439369150_15u
*******
.subckt 1510_74439370047_4.7u 1 2
Rp 1 2 4296
Cp 1 2 22.242p
Rs 1 N3 0.0031
L1 N3 2 4.217u
.ends 1510_74439370047_4.7u
*******
.subckt 1510_74439370068_6.8u 1 2
Rp 1 2 5066
Cp 1 2 21.801p
Rs 1 N3 0.0041
L1 N3 2 6.111u
.ends 1510_74439370068_6.8u
*******
.subckt 1510_74439370082_8.2u 1 2
Rp 1 2 6284
Cp 1 2 25.54p
Rs 1 N3 0.0055
L1 N3 2 8.328u
.ends 1510_74439370082_8.2u
*******
.subckt 1510_74439370100_10u 1 2
Rp 1 2 5244
Cp 1 2 29.045p
Rs 1 N3 0.0064
L1 N3 2 10.4u
.ends 1510_74439370100_10u
*******
.subckt 1510_74439370150_15u 1 2
Rp 1 2 7827
Cp 1 2 24.013p
Rs 1 N3 0.0105
L1 N3 2 15.895u
.ends 1510_74439370150_15u
*******
.subckt 1510_74439370220_22u 1 2
Rp 1 2 8204
Cp 1 2 26.195p
Rs 1 N3 0.0125
L1 N3 2 20.695u
.ends 1510_74439370220_22u
*******
.subckt 1510_74439370330_33u 1 2
Rp 1 2 10776
Cp 1 2 27.127p
Rs 1 N3 0.018
L1 N3 2 31.904u
.ends 1510_74439370330_33u
*******
.subckt 6030_744393440015_0.15u 1 2
Rp 1 2 306.09
Cp 1 2 4.722p
Rs 1 N3 0.00124
L1 N3 2 0.147u
.ends 6030_744393440015_0.15u
*******
.subckt 6030_744393440018_0.18u 1 2
Rp 1 2 393.041
Cp 1 2 5.062p
Rs 1 N3 0.00132
L1 N3 2 0.176u
.ends 6030_744393440018_0.18u
*******
.subckt 6030_744393440033_0.33u 1 2
Rp 1 2 683.781
Cp 1 2 6.324p
Rs 1 N3 0.0021
L1 N3 2 0.316u
.ends 6030_744393440033_0.33u
*******
.subckt 6030_744393440056_0.56u 1 2
Rp 1 2 876.79
Cp 1 2 7.515p
Rs 1 N3 0.0029
L1 N3 2 0.561u
.ends 6030_744393440056_0.56u
*******
.subckt 6030_74439344010_1u 1 2
Rp 1 2 1956
Cp 1 2 7.102p
Rs 1 N3 0.0055
L1 N3 2 1.008u
.ends 6030_74439344010_1u
*******
.subckt 6030_74439344012_1.2u 1 2
Rp 1 2 2178
Cp 1 2 8.182p
Rs 1 N3 0.0064
L1 N3 2 1.105u
.ends 6030_74439344012_1.2u
*******
.subckt 6030_74439344022_2.2u 1 2
Rp 1 2 2927
Cp 1 2 8.36p
Rs 1 N3 0.0105
L1 N3 2 2.182u
.ends 6030_74439344022_2.2u
*******
.subckt 6030_74439344033_3.3u 1 2
Rp 1 2 4970
Cp 1 2 7.979p
Rs 1 N3 0.0192
L1 N3 2 3.247u
.ends 6030_74439344033_3.3u
*******
.subckt 6030_74439344047_4.7u 1 2
Rp 1 2 7211
Cp 1 2 7.002p
Rs 1 N3 0.031
L1 N3 2 4.676u
.ends 6030_74439344047_4.7u
*******
.subckt 6060_74439346010_1u 1 2
Rp 1 2 1210
Cp 1 2 6.845p
Rs 1 N3 0.00339
L1 N3 2 1.046u
.ends 6060_74439346010_1u
*******
.subckt 6060_74439346012_1.2u 1 2
Rp 1 2 1330
Cp 1 2 8.78p
Rs 1 N3 0.00365
L1 N3 2 1.158u
.ends 6060_74439346012_1.2u
*******
.subckt 6060_74439346015_1.5u 1 2
Rp 1 2 1396
Cp 1 2 9.359p
Rs 1 N3 0.0039
L1 N3 2 1.373u
.ends 6060_74439346015_1.5u
*******
.subckt 6060_74439346018_1.8u 1 2
Rp 1 2 1659
Cp 1 2 7.994p
Rs 1 N3 0.0047
L1 N3 2 1.806u
.ends 6060_74439346018_1.8u
*******
.subckt 6060_74439346022_2.2u 1 2
Rp 1 2 1877
Cp 1 2 8.362p
Rs 1 N3 0.00558
L1 N3 2 2.182u
.ends 6060_74439346022_2.2u
*******
.subckt 6060_74439346033_3.3u 1 2
Rp 1 2 2955
Cp 1 2 8.785p
Rs 1 N3 0.01083
L1 N3 2 2.95u
.ends 6060_74439346033_3.3u
*******
.subckt 6060_74439346047_4.7u 1 2
Rp 1 2 4305
Cp 1 2 7.633p
Rs 1 N3 0.013
L1 N3 2 4.289u
.ends 6060_74439346047_4.7u
*******
.subckt 6060_74439346056_5.6u 1 2
Rp 1 2 5112
Cp 1 2 7.79p
Rs 1 N3 0.015
L1 N3 2 5.311u
.ends 6060_74439346056_5.6u
*******
.subckt 6060_74439346068_6.8u 1 2
Rp 1 2 5867
Cp 1 2 7.976p
Rs 1 N3 0.0176
L1 N3 2 6.553u
.ends 6060_74439346068_6.8u
*******
.subckt 6060_74439346082_8.2u 1 2
Rp 1 2 6820
Cp 1 2 8.668p
Rs 1 N3 0.023
L1 N3 2 7.855u
.ends 6060_74439346082_8.2u
*******
.subckt 6060_74439346100_10u 1 2
Rp 1 2 9786
Cp 1 2 8.192p
Rs 1 N3 0.0265
L1 N3 2 9.539u
.ends 6060_74439346100_10u
*******
.subckt 6060_74439346150_15u 1 2
Rp 1 2 11178
Cp 1 2 8.829p
Rs 1 N3 0.042
L1 N3 2 15.089u
.ends 6060_74439346150_15u
*******
.subckt 8080_744393580068_0.68u 1 2
Rp 1 2 1027
Cp 1 2 9.182p
Rs 1 N3 0.00141
L1 N3 2 0.71u
.ends 8080_744393580068_0.68u
*******
.subckt 8080_74439358010_1u 1 2
Rp 1 2 1445
Cp 1 2 8.916p
Rs 1 N3 0.0021
L1 N3 2 1.014u
.ends 8080_74439358010_1u
*******
.subckt 8080_74439358015_1.5u 1 2
Rp 1 2 1599
Cp 1 2 11.49p
Rs 1 N3 0.00291
L1 N3 2 1.588u
.ends 8080_74439358015_1.5u
*******
.subckt 8080_74439358022_2.2u 1 2
Rp 1 2 2282
Cp 1 2 10.434p
Rs 1 N3 0.0037
L1 N3 2 2.209u
.ends 8080_74439358022_2.2u
*******
.subckt 8080_74439358047_4.7u 1 2
Rp 1 2 4439
Cp 1 2 10.924p
Rs 1 N3 0.00865
L1 N3 2 4.785u
.ends 8080_74439358047_4.7u
*******
.subckt 8080_74439358068_6.8u 1 2
Rp 1 2 6545
Cp 1 2 7.924p
Rs 1 N3 0.013
L1 N3 2 6.596u
.ends 8080_74439358068_6.8u
*******
.subckt 8080_74439358100_10u 1 2
Rp 1 2 8417
Cp 1 2 8.116p
Rs 1 N3 0.019
L1 N3 2 10.282u
.ends 8080_74439358100_10u
*******
.subckt 8080_74439358150_15u 1 2
Rp 1 2 8485
Cp 1 2 11.885p
Rs 1 N3 0.025
L1 N3 2 14.163u
.ends 8080_74439358150_15u
*******
.subckt 4020_744393230022_0.22u 1 2
Rp 1 2 500
Cp 1 2 4.1p
Rs 1 N3 0.00305
L1 N3 2 0.231u
.ends 4020_744393230022_0.22u
*******
.subckt 4020_744393230047_0.47u 1 2
Rp 1 2 560.457
Cp 1 2 5.571p
Rs 1 N3 0.00525
L1 N3 2 0.47u
.ends 4020_744393230047_0.47u
*******
.subckt 4020_744393230056_0.56u 1 2
Rp 1 2 1264
Cp 1 2 6.009p
Rs 1 N3 0.0063
L1 N3 2 0.54u
.ends 4020_744393230056_0.56u
*******
.subckt 4020_744393230068_0.68u 1 2
Rp 1 2 1050
Cp 1 2 6.38p
Rs 1 N3 0.0066
L1 N3 2 0.63u
.ends 4020_744393230068_0.68u
*******
.subckt 4020_744393230082_0.82u 1 2
Rp 1 2 1325
Cp 1 2 6.414p
Rs 1 N3 0.0093
L1 N3 2 0.81u
.ends 4020_744393230082_0.82u
*******
.subckt 4020_74439323010_1u 1 2
Rp 1 2 1442
Cp 1 2 7.529p
Rs 1 N3 0.0107
L1 N3 2 1.03u
.ends 4020_74439323010_1u
*******
.subckt 4020_74439323012_1.2u 1 2
Rp 1 2 1678
Cp 1 2 7.325p
Rs 1 N3 0.0125
L1 N3 2 1.17u
.ends 4020_74439323012_1.2u
*******
.subckt 4020_74439323015_1.5u 1 2
Rp 1 2 2102
Cp 1 2 6.133p
Rs 1 N3 0.0163
L1 N3 2 1.44u
.ends 4020_74439323015_1.5u
*******
.subckt 4020_74439323022_2.2u 1 2
Rp 1 2 3075
Cp 1 2 8.237p
Rs 1 N3 0.0202
L1 N3 2 2.25u
.ends 4020_74439323022_2.2u
*******
.subckt 4030_744393240047_0.47u 1 2
Rp 1 2 707.603
Cp 1 2 5.023p
Rs 1 N3 0.0039
L1 N3 2 0.444u
.ends 4030_744393240047_0.47u
*******
.subckt 4030_744393240064_0.64u 1 2
Rp 1 2 1004
Cp 1 2 5.533p
Rs 1 N3 0.0048
L1 N3 2 0.591u
.ends 4030_744393240064_0.64u
*******
.subckt 4030_744393240090_0.90u 1 2
Rp 1 2 1043
Cp 1 2 7.898p
Rs 1 N3 0.0061
L1 N3 2 0.84u
.ends 4030_744393240090_0.90u
*******
.subckt 4030_74439324010_1u 1 2
Rp 1 2 1294
Cp 1 2 7.665p
Rs 1 N3 0.0087
L1 N3 2 0.65u
.ends 4030_74439324010_1u
*******
.subckt 4030_74439324012_1.2u 1 2
Rp 1 2 1507
Cp 1 2 7.672p
Rs 1 N3 0.0089
L1 N3 2 1.19u
.ends 4030_74439324012_1.2u
*******
.subckt 4030_74439324015_1.5u 1 2
Rp 1 2 1631
Cp 1 2 6.572p
Rs 1 N3 0.0101
L1 N3 2 1.37u
.ends 4030_74439324015_1.5u
*******
.subckt 4030_74439324022_2.2u 1 2
Rp 1 2 2709
Cp 1 2 7.314p
Rs 1 N3 0.0166
L1 N3 2 2.12u
.ends 4030_74439324022_2.2u
*******
.subckt 4030_74439324033_3.3u 1 2
Rp 1 2 2911
Cp 1 2 8.896p
Rs 1 N3 0.0202
L1 N3 2 3.26u
.ends 4030_74439324033_3.3u
*******
.subckt 4030_74439324047_4.7u 1 2
Rp 1 2 6900
Cp 1 2 7.185p
Rs 1 N3 0.0313
L1 N3 2 4.49u
.ends 4030_74439324047_4.7u
*******
.subckt 4040_74439325033_3.3u 1 2
Rp 1 2 2925
Cp 1 2 8.544p
Rs 1 N3 0.0204
L1 N3 2 3.217u
.ends 4040_74439325033_3.3u
*******
.subckt 4040_74439325047_4.7u 1 2
Rp 1 2 2552
Cp 1 2 9.462p
Rs 1 N3 0.0265
L1 N3 2 4.966u
.ends 4040_74439325047_4.7u
*******
.subckt 4040_74439325056_5.6u 1 2
Rp 1 2 6407
Cp 1 2 8.287p
Rs 1 N3 0.0342
L1 N3 2 5.719u
.ends 4040_74439325056_5.6u
*******
.subckt 4040_74439325068_6.8u 1 2
Rp 1 2 10604
Cp 1 2 6.978p
Rs 1 N3 0.0423
L1 N3 2 6.707u
.ends 4040_74439325068_6.8u
*******
.subckt 5020_744393330016_0.16u 1 2
Rp 1 2 332.836
Cp 1 2 4.771p
Rs 1 N3 0.0022
L1 N3 2 0.148u
.ends 5020_744393330016_0.16u
*******
.subckt 5020_744393330033_0.33u 1 2
Rp 1 2 546.947
Cp 1 2 7.165p
Rs 1 N3 0.003
L1 N3 2 0.332u
.ends 5020_744393330033_0.33u
*******
.subckt 5020_744393330056_0.56u 1 2
Rp 1 2 849.046
Cp 1 2 5.993p
Rs 1 N3 0.0052
L1 N3 2 0.536u
.ends 5020_744393330056_0.56u
*******
.subckt 5020_744393330068_0.68u 1 2
Rp 1 2 1181
Cp 1 2 6.54p
Rs 1 N3 0.0067
L1 N3 2 0.72u
.ends 5020_744393330068_0.68u
*******
.subckt 5020_74439333010_1u 1 2
Rp 1 2 950
Cp 1 2 9.636p
Rs 1 N3 0.0095
L1 N3 2 0.97u
.ends 5020_74439333010_1u
*******
.subckt 5020_74439333012_1.2u 1 2
Rp 1 2 1708
Cp 1 2 8.409p
Rs 1 N3 0.0108
L1 N3 2 1.25u
.ends 5020_74439333012_1.2u
*******
.subckt 5030_744393340033_0.33u 1 2
Rp 1 2 574.378
Cp 1 2 7.026p
Rs 1 N3 0.00301
L1 N3 2 0.328238u
.ends 5030_744393340033_0.33u
*******
.subckt 5030_744393340056_0.56u 1 2
Rp 1 2 836.509
Cp 1 2 8.126p
Rs 1 N3 0.00399
L1 N3 2 0.546969u
.ends 5030_744393340056_0.56u
*******
.subckt 5030_744393340068_0.68u 1 2
Rp 1 2 613.431
Cp 1 2 9.363p
Rs 1 N3 0.00409
L1 N3 2 0.691759u
.ends 5030_744393340068_0.68u
*******
.subckt 5030_74439334010_1u 1 2
Rp 1 2 810.15
Cp 1 2 10.541p
Rs 1 N3 0.0063
L1 N3 2 0.66854u
.ends 5030_74439334010_1u
*******
.subckt 5030_74439334012_1.2u 1 2
Rp 1 2 1486
Cp 1 2 9.582p
Rs 1 N3 0.0066
L1 N3 2 1.219u
.ends 5030_74439334012_1.2u
*******
.subckt 5030_74439334015_1.5u 1 2
Rp 1 2 1932
Cp 1 2 8.871p
Rs 1 N3 0.008
L1 N3 2 1.614u
.ends 5030_74439334015_1.5u
*******
.subckt 5030_74439334022_2.2u 1 2
Rp 1 2 2762
Cp 1 2 9.83p
Rs 1 N3 0.0113
L1 N3 2 2.13u
.ends 5030_74439334022_2.2u
*******
.subckt 5030_74439334033_3.3u 1 2
Rp 1 2 2140
Cp 1 2 11.045p
Rs 1 N3 0.0163
L1 N3 2 3.496u
.ends 5030_74439334033_3.3u
*******
.subckt 5030_74439334047_4.7u 1 2
Rp 1 2 3991
Cp 1 2 10.549p
Rs 1 N3 0.0229
L1 N3 2 4.943u
.ends 5030_74439334047_4.7u
*******
.subckt 5050_744393305056_5.6u 1 2
Rp 1 2 3527
Cp 1 2 9.72p
Rs 1 N3 0.0218
L1 N3 2 5.702u
.ends 5050_744393305056_5.6u
*******
.subckt 5050_744393305068_6.8u 1 2
Rp 1 2 9422
Cp 1 2 11.47p
Rs 1 N3 0.0237
L1 N3 2 6.846u
.ends 5050_744393305068_6.8u
*******
.subckt 5050_744393305082_8.2u 1 2
Rp 1 2 11476
Cp 1 2 10.965p
Rs 1 N3 0.0293
L1 N3 2 8.338u
.ends 5050_744393305082_8.2u
*******
.subckt 5050_744393305100_10u 1 2
Rp 1 2 4502
Cp 1 2 12.201p
Rs 1 N3 0.0354
L1 N3 2 10.647u
.ends 5050_744393305100_10u
*******
.subckt 5050_744393305150_15u 1 2
Rp 1 2 17051
Cp 1 2 10.749p
Rs 1 N3 0.0568
L1 N3 2 16.504u
.ends 5050_744393305150_15u
*******
.subckt 5050_744393305220_22u 1 2
Rp 1 2 19323
Cp 1 2 11.699p
Rs 1 N3 0.075
L1 N3 2 22.094u
.ends 5050_744393305220_22u
*******
.subckt 7030_74439384010_1u 1 2
Rp 1 2 1583
Cp 1 2 11.684p
Rs 1 N3 0.0039
L1 N3 2 0.9456u
.ends 7030_74439384010_1u
*******
.subckt 7030_74439384012_1.2u 1 2
Rp 1 2 841
Cp 1 2 14.189p
Rs 1 N3 0.0042
L1 N3 2 1.157u
.ends 7030_74439384012_1.2u
*******
.subckt 7030_74439384015_1.5u 1 2
Rp 1 2 1847
Cp 1 2 11.892p
Rs 1 N3 0.0051
L1 N3 2 1.393u
.ends 7030_74439384015_1.5u
*******
.subckt 7030_74439384022_2.2u 1 2
Rp 1 2 2530
Cp 1 2 14.021p
Rs 1 N3 0.0079
L1 N3 2 2.223u
.ends 7030_74439384022_2.2u
*******
.subckt 7030_74439384033_3.3u 1 2
Rp 1 2 3242
Cp 1 2 12.561p
Rs 1 N3 0.0144
L1 N3 2 3.171u
.ends 7030_74439384033_3.3u
*******
.subckt 7030_74439384047_4.7u 1 2
Rp 1 2 5033
Cp 1 2 13.362p
Rs 1 N3 0.0198
L1 N3 2 5.149u
.ends 7030_74439384047_4.7u
*******
.subckt 7070_74439387033_3.3u 1 2
Rp 1 2 2426
Cp 1 2 14.688p
Rs 1 N3 0.0064
L1 N3 2 3.212u
.ends 7070_74439387033_3.3u
*******
.subckt 7070_74439387047_4.7u 1 2
Rp 1 2 3245
Cp 1 2 13.478p
Rs 1 N3 0.0092
L1 N3 2 4.617u
.ends 7070_74439387047_4.7u
*******
.subckt 7070_74439387056_5.6u 1 2
Rp 1 2 2248
Cp 1 2 18.924p
Rs 1 N3 0.0124
L1 N3 2 5.67u
.ends 7070_74439387056_5.6u
*******
.subckt 7070_74439387068_6.8u 1 2
Rp 1 2 2887
Cp 1 2 15.001p
Rs 1 N3 0.0124
L1 N3 2 6.749u
.ends 7070_74439387068_6.8u
*******
.subckt 7070_74439387082_8.2u 1 2
Rp 1 2 3645
Cp 1 2 16.219p
Rs 1 N3 0.0145
L1 N3 2 8.537u
.ends 7070_74439387082_8.2u
*******
.subckt 7070_74439387100_10u 1 2
Rp 1 2 4865
Cp 1 2 14.504p
Rs 1 N3 0.019
L1 N3 2 9.866u
.ends 7070_74439387100_10u
*******