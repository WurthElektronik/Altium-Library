**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ASLL
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         5/31/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 865060140001_22uF 1 2
Rser 1 3 1.95778285719
Lser 2 4 1.32310492E-09
C1 3 4 0.000022
Rpar 3 4 2100000
.ends 865060140001_22uF
*******
.subckt 865060140002_33uF 1 2
Rser 1 3 1.39
Lser 2 4 9.94648012E-10
C1 3 4 0.000033
Rpar 3 4 2100000
.ends 865060140002_33uF
*******
.subckt 865060142003_47uF 1 2
Rser 1 3 0.93
Lser 2 4 0.000000002268
C1 3 4 0.000047
Rpar 3 4 2100000
.ends 865060142003_47uF
*******
.subckt 865060143004_100uF 1 2
Rser 1 3 0.52
Lser 2 4 0.000000002445
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865060143004_100uF
*******
.subckt 865060143005_150uF 1 2
Rser 1 3 0.43
Lser 2 4 0.000000002568
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865060143005_150uF
*******
.subckt 865060145006_220uF 1 2
Rser 1 3 0.215
Lser 2 4 4.89349029708004E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865060145006_220uF
*******
.subckt 865060153007_330uF 1 2
Rser 1 3 0.115
Lser 2 4 6.07922445196185E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865060153007_330uF
*******
.subckt 865060153008_470uF 1 2
Rser 1 3 0.114
Lser 2 4 6.33636829390827E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865060153008_470uF
*******
.subckt 865060153009_680uF 1 2
Rser 1 3 0.102
Lser 2 4 6.30794647678417E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865060153009_680uF
*******
.subckt 865060153010_1mF 1 2
Rser 1 3 0.15277116107
Lser 2 4 6.41430176E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 865060153010_1mF
*******
.subckt 865060157011_1.5mF 1 2
Rser 1 3 0.071
Lser 2 4 6.62915805201144E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 865060157011_1.5mF
*******
.subckt 865060162012_3.3mF 1 2
Rser 1 3 0.0883426572544
Lser 2 4 1.1533778839E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 865060162012_3.3mF
*******
.subckt 865060163013_6.8mF 1 2
Rser 1 3 0.0491759976628
Lser 2 4 1.4371157676E-08
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 865060163013_6.8mF
*******
.subckt 865060240001_22uF 1 2
Rser 1 3 1.97248561552
Lser 2 4 1.225987906E-09
C1 3 4 0.000022
Rpar 3 4 3333333.33333333
.ends 865060240001_22uF
*******
.subckt 865060242002_33uF 1 2
Rser 1 3 0.85
Lser 2 4 1.749069264E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865060242002_33uF
*******
.subckt 865060243003_47uF 1 2
Rser 1 3 0.413
Lser 2 4 1.90914369178307E-08
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865060243003_47uF
*******
.subckt 865060243004_100uF 1 2
Rser 1 3 0.48
Lser 2 4 0.000000002516
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865060243004_100uF
*******
.subckt 865060243005_150uF 1 2
Rser 1 3 0.49
Lser 2 4 0.000000002554
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865060243005_150uF
*******
.subckt 865060245006_220uF 1 2
Rser 1 3 0.377
Lser 2 4 2.807249688E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865060245006_220uF
*******
.subckt 865060253007_330uF 1 2
Rser 1 3 0.122
Lser 2 4 5.88662119916188E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865060253007_330uF
*******
.subckt 865060253008_470uF 1 2
Rser 1 3 0.104
Lser 2 4 6.47919311195411E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865060253008_470uF
*******
.subckt 865060257009_680uF 1 2
Rser 1 3 0.068
Lser 2 4 7.47892860793178E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865060257009_680uF
*******
.subckt 865060257010_1mF 1 2
Rser 1 3 0.134172089212
Lser 2 4 7.553834187E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 865060257010_1mF
*******
.subckt 865060262011_2.2mF 1 2
Rser 1 3 0.0849933988011
Lser 2 4 1.3636764258E-08
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 865060262011_2.2mF
*******
.subckt 865060263012_4.7mF 1 2
Rser 1 3 0.0453775892498
Lser 2 4 1.7398862797E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 865060263012_4.7mF
*******
.subckt 865060340001_10uF 1 2
Rser 1 3 1.82554735976
Lser 2 4 2.122293627E-09
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 865060340001_10uF
*******
.subckt 865060342002_22uF 1 2
Rser 1 3 1.20935467322
Lser 2 4 1.666028416E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865060342002_22uF
*******
.subckt 865060343003_33uF 1 2
Rser 1 3 0.5
Lser 2 4 0.000000002457
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865060343003_33uF
*******
.subckt 865060343004_47uF 1 2
Rser 1 3 0.432
Lser 2 4 0.000000002917
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865060343004_47uF
*******
.subckt 865060343005_100uF 1 2
Rser 1 3 0.339
Lser 2 4 1.92595385133346E-08
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865060343005_100uF
*******
.subckt 865060345006_150uF 1 2
Rser 1 3 0.261
Lser 2 4 4.17226894584708E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865060345006_150uF
*******
.subckt 865060345007_220uF 1 2
Rser 1 3 0.255
Lser 2 4 2.0004545428038E-08
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865060345007_220uF
*******
.subckt 865060353008_330uF 1 2
Rser 1 3 0.114
Lser 2 4 7.04229949303687E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865060353008_330uF
*******
.subckt 865060353009_470uF 1 2
Rser 1 3 0.106
Lser 2 4 6.11214672792288E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865060353009_470uF
*******
.subckt 865060357010_680uF 1 2
Rser 1 3 0.076
Lser 2 4 7.54382183012106E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865060357010_680uF
*******
.subckt 865060362011_1.5mF 1 2
Rser 1 3 0.0746402783307
Lser 2 4 1.1233002286E-08
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 865060362011_1.5mF
*******
.subckt 865060363012_3.3mF 1 2
Rser 1 3 0.0506090430045
Lser 2 4 1.7281079821E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 865060363012_3.3mF
*******
.subckt 865060440001_10uF 1 2
Rser 1 3 1.81968584275
Lser 2 4 1.435032181E-09
C1 3 4 0.00001
Rpar 3 4 8333333.33333333
.ends 865060440001_10uF
*******
.subckt 865060442002_22uF 1 2
Rser 1 3 0.87731
Lser 2 4 1.829921963E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865060442002_22uF
*******
.subckt 865060443003_33uF 1 2
Rser 1 3 0.425
Lser 2 4 0.000000002581
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865060443003_33uF
*******
.subckt 865060443004_47uF 1 2
Rser 1 3 0.49577
Lser 2 4 2.561764526E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865060443004_47uF
*******
.subckt 865060445005_100uF 1 2
Rser 1 3 0.248
Lser 2 4 4.65325272922483E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865060445005_100uF
*******
.subckt 865060453006_150uF 1 2
Rser 1 3 0.131
Lser 2 4 5.32075249490287E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865060453006_150uF
*******
.subckt 865060453007_220uF 1 2
Rser 1 3 0.115
Lser 2 4 6.11819272741701E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865060453007_220uF
*******
.subckt 865060453008_330uF 1 2
Rser 1 3 0.104
Lser 2 4 6.41491656365575E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865060453008_330uF
*******
.subckt 865060457009_470uF 1 2
Rser 1 3 0.075
Lser 2 4 6.99799142847963E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865060457009_470uF
*******
.subckt 865060462010_1mF 1 2
Rser 1 3 0.0680864476895
Lser 2 4 1.0639515132E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 865060462010_1mF
*******
.subckt 865060463011_2.2mF 1 2
Rser 1 3 0.0456127811975
Lser 2 4 1.3570666657E-08
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 865060463011_2.2mF
*******
.subckt 865060540001_4.7uF 1 2
Rser 1 3 1.51
Lser 2 4 0.000000000908767
C1 3 4 0.0000047
Rpar 3 4 11666666.6666667
.ends 865060540001_4.7uF
*******
.subckt 865060542002_10uF 1 2
Rser 1 3 0.8
Lser 2 4 1.753067519E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865060542002_10uF
*******
.subckt 865060543003_22uF 1 2
Rser 1 3 0.46358
Lser 2 4 2.631136726E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 865060543003_22uF
*******
.subckt 865060543004_33uF 1 2
Rser 1 3 0.396
Lser 2 4 1.8322629471383E-08
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865060543004_33uF
*******
.subckt 865060543005_47uF 1 2
Rser 1 3 0.32
Lser 2 4 0.000000002746
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865060543005_47uF
*******
.subckt 865060553006_100uF 1 2
Rser 1 3 0.104
Lser 2 4 5.87152525559351E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865060553006_100uF
*******
.subckt 865060553007_150uF 1 2
Rser 1 3 0.108
Lser 2 4 6.32536831819924E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865060553007_150uF
*******
.subckt 865060557008_220uF 1 2
Rser 1 3 0.101928277741
Lser 2 4 8.987682735E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865060557008_220uF
*******
.subckt 865060562009_470uF 1 2
Rser 1 3 0.0614283665816
Lser 2 4 1.089209523E-08
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865060562009_470uF
*******
.subckt 865060562010_680uF 1 2
Rser 1 3 0.0623680408299
Lser 2 4 1.0309509399E-08
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865060562010_680uF
*******
.subckt 865060563011_1mF 1 2
Rser 1 3 0.07287
Lser 2 4 3.7385992735E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 865060563011_1mF
*******
.subckt 865060563012_1.5mF 1 2
Rser 1 3 0.0421315277337
Lser 2 4 1.3525660889E-08
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 865060563012_1.5mF
*******
.subckt 865060640001_1uF 1 2
Rser 1 3 2.2635885173
Lser 2 4 1.360271975E-09
C1 3 4 0.000001
Rpar 3 4 16666666.6666667
.ends 865060640001_1uF
*******
.subckt 865060640002_2.2uF 1 2
Rser 1 3 2.3327154948
Lser 2 4 1.352818032E-09
C1 3 4 0.0000022
Rpar 3 4 16666666.6666667
.ends 865060640002_2.2uF
*******
.subckt 865060640003_3.3uF 1 2
Rser 1 3 2.28875666379
Lser 2 4 1.338582645E-09
C1 3 4 0.0000033
Rpar 3 4 16666666.6666667
.ends 865060640003_3.3uF
*******
.subckt 865060642004_4.7uF 1 2
Rser 1 3 1.4
Lser 2 4 0.000000001219
C1 3 4 0.0000047
Rpar 3 4 16666666.6666667
.ends 865060642004_4.7uF
*******
.subckt 865060643005_10uF 1 2
Rser 1 3 0.86
Lser 2 4 0.000000002536
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865060643005_10uF
*******
.subckt 865060643006_22uF 1 2
Rser 1 3 0.885
Lser 2 4 0.000000002678
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865060643006_22uF
*******
.subckt 865060645007_33uF 1 2
Rser 1 3 0.59
Lser 2 4 0.000000002434
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865060645007_33uF
*******
.subckt 865060645008_47uF 1 2
Rser 1 3 0.47
Lser 2 4 0.000000002471
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865060645008_47uF
*******
.subckt 865060653009_68uF 1 2
Rser 1 3 0.235
Lser 2 4 4.89808349206542E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 865060653009_68uF
*******
.subckt 865060653010_100uF 1 2
Rser 1 3 0.196
Lser 2 4 5.50548674447443E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865060653010_100uF
*******
.subckt 865060657011_150uF 1 2
Rser 1 3 0.14
Lser 2 4 6.4296689103223E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865060657011_150uF
*******
.subckt 865060657012_220uF 1 2
Rser 1 3 0.152
Lser 2 4 1.32310492E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865060657012_220uF
*******
.subckt 865060663013_470uF 1 2
Rser 1 3 0.0689885274662
Lser 2 4 6.625564537E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865060663013_470uF
*******
.subckt 865060663014_680uF 1 2
Rser 1 3 0.0676767846067
Lser 2 4 1.4060641893E-08
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865060663014_680uF
*******
.subckt 865060663015_1mF 1 2
Rser 1 3 0.0672430678769
Lser 2 4 1.3729957932E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 865060663015_1mF
*******
.subckt 865060742001_4.7uF 1 2
Rser 1 3 2.19830173265
Lser 2 4 1.510333447E-09
C1 3 4 0.0000047
Rpar 3 4 21000000
.ends 865060742001_4.7uF
*******
.subckt 865060743002_10uF 1 2
Rser 1 3 1.15438062397
Lser 2 4 2.120138712E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865060743002_10uF
*******
.subckt 865060745003_22uF 1 2
Rser 1 3 0.629
Lser 2 4 2.584346505E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865060745003_22uF
*******
.subckt 865060753004_33uF 1 2
Rser 1 3 0.44486
Lser 2 4 3.333290236E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865060753004_33uF
*******
.subckt 865060753005_47uF 1 2
Rser 1 3 0.295
Lser 2 4 3.477908007E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865060753005_47uF
*******
.subckt 865060757006_68uF 1 2
Rser 1 3 0.25696
Lser 2 4 4.629373515E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 865060757006_68uF
*******
.subckt 865060757007_100uF 1 2
Rser 1 3 0.22141
Lser 2 4 6.564382958E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865060757007_100uF
*******
.subckt 865060762008_150uF 1 2
Rser 1 3 0.14542
Lser 2 4 6.42301006E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865060762008_150uF
*******
.subckt 865060762009_220uF 1 2
Rser 1 3 0.18803
Lser 2 4 6.625564537E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865060762009_220uF
*******
.subckt 865060763010_470uF 1 2
Rser 1 3 0.0715
Lser 2 4 1.2835672547E-08
C1 3 4 0.00047
Rpar 3 4 212765.957446808
.ends 865060763010_470uF
*******
.subckt 865060845002_10uF 1 2
Rser 1 3 1.23100255905
Lser 2 4 2.141910579E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865060845002_10uF
*******
.subckt 865060853003_22uF 1 2
Rser 1 3 0.994
Lser 2 4 2.860638601E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865060853003_22uF
*******
.subckt 865060857004_33uF 1 2
Rser 1 3 0.83111
Lser 2 4 3.664633085E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865060857004_33uF
*******
.subckt 865060857005_47uF 1 2
Rser 1 3 0.83611
Lser 2 4 5.230622691E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865060857005_47uF
*******
.subckt 865060862006_68uF 1 2
Rser 1 3 0.377
Lser 2 4 5.633545651E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 865060862006_68uF
*******
.subckt 865061457001_3.3uF 1 2
Rser 1 3 0.98034
Lser 2 4 4.014064484E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 865061457001_3.3uF
*******
.subckt 865061462002_4.7uF 1 2
Rser 1 3 0.8763
Lser 2 4 5.53708126E-09
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 865061462002_4.7uF
*******
.subckt 865061462003_6.8uF 1 2
Rser 1 3 0.88125
Lser 2 4 5.106986815E-09
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 865061462003_6.8uF
*******
.subckt 865061462004_10uF 1 2
Rser 1 3 1.05493385794
Lser 2 4 1.1650705766E-08
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865061462004_10uF
*******
.subckt 865061463005_15uF 1 2
Rser 1 3 0.57464
Lser 2 4 6.64629781E-09
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends 865061463005_15uF
*******
