**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT Power Inductor
* Matchcode:             WE-PD2A
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         2021/06/09
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1054_784776047_4.7u 1 2
Rp 1 2 7013
Cp 1 2 3.36986p
Rs 1 N3 0.012
L1 N3 2 3.589u
.ends 1054_784776047_4.7u
*******
.subckt 1054_784776056_5.6u 1 2
Rp 1 2 8735
Cp 1 2 3.21304p
Rs 1 N3 0.015
L1 N3 2 4.384u
.ends 1054_784776056_5.6u
*******
.subckt 1054_784776068_6.8u 1 2
Rp 1 2 10473
Cp 1 2 4.92116p
Rs 1 N3 0.016
L1 N3 2 5.426u
.ends 1054_784776068_6.8u
*******
.subckt 1054_784776082_8.2u 1 2
Rp 1 2 13497
Cp 1 2 4.69346p
Rs 1 N3 0.02
L1 N3 2 7.272u
.ends 1054_784776082_8.2u
*******
.subckt 1054_78477610_10u 1 2
Rp 1 2 13035
Cp 1 2 3.80778p
Rs 1 N3 0.028
L1 N3 2 8.658u
.ends 1054_78477610_10u
*******
.subckt 1054_784776112_12u 1 2
Rp 1 2 19542
Cp 1 2 3.77p
Rs 1 N3 0.033
L1 N3 2 9.935u
.ends 1054_784776112_12u
*******
.subckt 1054_784776115_15u 1 2
Rp 1 2 20035
Cp 1 2 5.34314p
Rs 1 N3 0.034
L1 N3 2 12.552u
.ends 1054_784776115_15u
*******
.subckt 1054_784776118_18u 1 2
Rp 1 2 23601
Cp 1 2 5.93414p
Rs 1 N3 0.043
L1 N3 2 15.658u
.ends 1054_784776118_18u
*******
.subckt 1054_784776122_22u 1 2
Rp 1 2 25733
Cp 1 2 5.51588p
Rs 1 N3 0.051
L1 N3 2 18.451u
.ends 1054_784776122_22u
*******
.subckt 1054_784776127_27u 1 2
Rp 1 2 32972
Cp 1 2 6.03448p
Rs 1 N3 0.063
L1 N3 2 12.266u
.ends 1054_784776127_27u
*******
.subckt 1054_784776133_33u 1 2
Rp 1 2 31667
Cp 1 2 5.84886p
Rs 1 N3 0.083
L1 N3 2 29.335u
.ends 1054_784776133_33u
*******
.subckt 1054_784776139_39u 1 2
Rp 1 2 42128
Cp 1 2 6.33974p
Rs 1 N3 0.098
L1 N3 2 33.497u
.ends 1054_784776139_39u
*******
.subckt 1054_784776147_47u 1 2
Rp 1 2 48128
Cp 1 2 7.16597p
Rs 1 N3 0.095
L1 N3 2 37.549u
.ends 1054_784776147_47u
*******
.subckt 1054_784776156_56u 1 2
Rp 1 2 56398
Cp 1 2 6.50986p
Rs 1 N3 0.112
L1 N3 2 46.375u
.ends 1054_784776156_56u
*******
.subckt 1054_784776168_68u 1 2
Rp 1 2 48869
Cp 1 2 6.13886p
Rs 1 N3 0.138
L1 N3 2 54.849u
.ends 1054_784776168_68u
*******
.subckt 1054_784776182_82u 1 2
Rp 1 2 67716
Cp 1 2 7.76986p
Rs 1 N3 0.15
L1 N3 2 64.367u
.ends 1054_784776182_82u
*******
.subckt 1054_78477620_100u 1 2
Rp 1 2 60028
Cp 1 2 6.84462p
Rs 1 N3 0.2
L1 N3 2 83.124u
.ends 1054_78477620_100u
*******
.subckt 1054_784776212_120u 1 2
Rp 1 2 85667
Cp 1 2 7.64003p
Rs 1 N3 0.243
L1 N3 2 94.482u
.ends 1054_784776212_120u
*******
.subckt 1054_784776215_150u 1 2
Rp 1 2 102377
Cp 1 2 6.22604p
Rs 1 N3 0.3
L1 N3 2 132.75u
.ends 1054_784776215_150u
*******
.subckt 1054_784776218_180u 1 2
Rp 1 2 92907
Cp 1 2 6.5131p
Rs 1 N3 0.32
L1 N3 2 157.07u
.ends 1054_784776218_180u
*******
.subckt 1054_784776222_220u 1 2
Rp 1 2 93099
Cp 1 2 6.77668p
Rs 1 N3 0.451
L1 N3 2 186.036u
.ends 1054_784776222_220u
*******
.subckt 1054_784776227_270u 1 2
Rp 1 2 89759
Cp 1 2 7.93p
Rs 1 N3 0.5
L1 N3 2 212.716u
.ends 1054_784776227_270u
*******
.subckt 1054_784776233_330u 1 2
Rp 1 2 141012
Cp 1 2 6.8493p
Rs 1 N3 0.75
L1 N3 2 295.178u
.ends 1054_784776233_330u
*******
.subckt 1054_784776239_390u 1 2
Rp 1 2 149517
Cp 1 2 7.90624p
Rs 1 N3 0.794
L1 N3 2 329.891u
.ends 1054_784776239_390u
*******
.subckt 1054_784776247_470u 1 2
Rp 1 2 137510
Cp 1 2 7.32854p
Rs 1 N3 0.969
L1 N3 2 407.65u
.ends 1054_784776247_470u
*******
.subckt 4532_7847730_1u 1 2
Rp 1 2 4148
Cp 1 2 1.199p
Rs 1 N3 0.014
L1 N3 2 0.82036u
.ends 4532_7847730_1u
*******
.subckt 4532_784773018_1.8u 1 2
Rp 1 2 5754
Cp 1 2 1.5247p
Rs 1 N3 0.028
L1 N3 2 1.329u
.ends 4532_784773018_1.8u
*******
.subckt 4532_784773022_2.2u 1 2
Rp 1 2 6715
Cp 1 2 1.577p
Rs 1 N3 0.034
L1 N3 2 1.639u
.ends 4532_784773022_2.2u
*******
.subckt 4532_784773033_3.3u 1 2
Rp 1 2 10323
Cp 1 2 1.663p
Rs 1 N3 0.041
L1 N3 2 2.837u
.ends 4532_784773033_3.3u
*******
.subckt 4532_784773039_3.9u 1 2
Rp 1 2 10621
Cp 1 2 1.631p
Rs 1 N3 0.054
L1 N3 2 3.049u
.ends 4532_784773039_3.9u
*******
.subckt 4532_784773047_4.7u 1 2
Rp 1 2 12896
Cp 1 2 1.656p
Rs 1 N3 0.059
L1 N3 2 4.008u
.ends 4532_784773047_4.7u
*******
.subckt 4532_784773056_5.6u 1 2
Rp 1 2 14249
Cp 1 2 1.67p
Rs 1 N3 0.069
L1 N3 2 4.467u
.ends 4532_784773056_5.6u
*******
.subckt 4532_784773068_6.8u 1 2
Rp 1 2 17041
Cp 1 2 1.774p
Rs 1 N3 0.076
L1 N3 2 5.832u
.ends 4532_784773068_6.8u
*******
.subckt 4532_784773082_8.2u 1 2
Rp 1 2 18807
Cp 1 2 2.082p
Rs 1 N3 0.116
L1 N3 2 7.123u
.ends 4532_784773082_8.2u
*******
.subckt 4532_78477310_10u 1 2
Rp 1 2 22283
Cp 1 2 1.951p
Rs 1 N3 0.118
L1 N3 2 8.484u
.ends 4532_78477310_10u
*******
.subckt 4532_784773112_12u 1 2
Rp 1 2 21994
Cp 1 2 1.954p
Rs 1 N3 0.156
L1 N3 2 8.487u
.ends 4532_784773112_12u
*******
.subckt 4532_784773115_15u 1 2
Rp 1 2 27492
Cp 1 2 2.136p
Rs 1 N3 0.204
L1 N3 2 12.605u
.ends 4532_784773115_15u
*******
.subckt 4532_784773118_18u 1 2
Rp 1 2 32281
Cp 1 2 2.023p
Rs 1 N3 0.225
L1 N3 2 15.888u
.ends 4532_784773118_18u
*******
.subckt 4532_784773122_22u 1 2
Rp 1 2 37300
Cp 1 2 2.165p
Rs 1 N3 0.261
L1 N3 2 18.765u
.ends 4532_784773122_22u
*******
.subckt 4532_784773127_27u 1 2
Rp 1 2 38285
Cp 1 2 2.094p
Rs 1 N3 0.328
L1 N3 2 21.785u
.ends 4532_784773127_27u
*******
.subckt 4532_784773133_33u 1 2
Rp 1 2 38224
Cp 1 2 2.087p
Rs 1 N3 0.37
L1 N3 2 21.829u
.ends 4532_784773133_33u
*******
.subckt 4532_784773139_39u 1 2
Rp 1 2 49291
Cp 1 2 9.889p
Rs 1 N3 0.418
L1 N3 2 24.645u
.ends 4532_784773139_39u
*******
.subckt 4532_784773147_47u 1 2
Rp 1 2 74067
Cp 1 2 2.231p
Rs 1 N3 0.523
L1 N3 2 40.081u
.ends 4532_784773147_47u
*******
.subckt 4532_784773156_56u 1 2
Rp 1 2 65219
Cp 1 2 2.383p
Rs 1 N3 0.714
L1 N3 2 48.363u
.ends 4532_784773156_56u
*******
.subckt 4532_784773168_68u 1 2
Rp 1 2 73900
Cp 1 2 2.431p
Rs 1 N3 0.754
L1 N3 2 67.063u
.ends 4532_784773168_68u
*******
.subckt 5848_784774003_0.33u 1 2
Rp 1 2 2639
Cp 1 2 1.009p
Rs 1 N3 0.006
L1 N3 2 0.275482u
.ends 5848_784774003_0.33u
*******
.subckt 5848_784774006_0.6u 1 2
Rp 1 2 3985
Cp 1 2 1.085p
Rs 1 N3 0.009
L1 N3 2 0.453226u
.ends 5848_784774006_0.6u
*******
.subckt 5848_784774022_2.2u 1 2
Rp 1 2 11653
Cp 1 2 2.969p
Rs 1 N3 0.026
L1 N3 2 1.943u
.ends 5848_784774022_2.2u
*******
.subckt 5848_784774027_2.7u 1 2
Rp 1 2 12943
Cp 1 2 3.278p
Rs 1 N3 0.032
L1 N3 2 2.396u
.ends 5848_784774027_2.7u
*******
.subckt 5848_784774033_3.3u 1 2
Rp 1 2 15188
Cp 1 2 3.369p
Rs 1 N3 0.042
L1 N3 2 2.942u
.ends 5848_784774033_3.3u
*******
.subckt 5848_784774047_4.7u 1 2
Rp 1 2 18558
Cp 1 2 3.497p
Rs 1 N3 0.056
L1 N3 2 4.074u
.ends 5848_784774047_4.7u
*******
.subckt 5848_784774068_6.8u 1 2
Rp 1 2 22018
Cp 1 2 3.263p
Rs 1 N3 0.071
L1 N3 2 5.258u
.ends 5848_784774068_6.8u
*******
.subckt 5848_78477410_10u 1 2
Rp 1 2 18212
Cp 1 2 2.667p
Rs 1 N3 0.078
L1 N3 2 8.486u
.ends 5848_78477410_10u
*******
.subckt 5848_784774112_12u 1 2
Rp 1 2 20530
Cp 1 2 2.69p
Rs 1 N3 0.082
L1 N3 2 9.635u
.ends 5848_784774112_12u
*******
.subckt 5848_784774115_15u 1 2
Rp 1 2 28976
Cp 1 2 2.836p
Rs 1 N3 0.089
L1 N3 2 13.236u
.ends 5848_784774115_15u
*******
.subckt 5848_784774118_18u 1 2
Rp 1 2 28884
Cp 1 2 2.86p
Rs 1 N3 0.104
L1 N3 2 15.413u
.ends 5848_784774118_18u
*******
.subckt 5848_784774122_22u 1 2
Rp 1 2 35680
Cp 1 2 2.97p
Rs 1 N3 0.109
L1 N3 2 18.8u
.ends 5848_784774122_22u
*******
.subckt 5848_784774127_27u 1 2
Rp 1 2 45599
Cp 1 2 3.334p
Rs 1 N3 0.133
L1 N3 2 24.478u
.ends 5848_784774127_27u
*******
.subckt 5848_784774133_33u 1 2
Rp 1 2 53466
Cp 1 2 3.138p
Rs 1 N3 0.15
L1 N3 2 31.073u
.ends 5848_784774133_33u
*******
.subckt 5848_784774139_39u 1 2
Rp 1 2 51434
Cp 1 2 2.866p
Rs 1 N3 0.215
L1 N3 2 34.953u
.ends 5848_784774139_39u
*******
.subckt 5848_784774147_47u 1 2
Rp 1 2 54986
Cp 1 2 3.003p
Rs 1 N3 0.26
L1 N3 2 39.885u
.ends 5848_784774147_47u
*******
.subckt 5848_784774156_56u 1 2
Rp 1 2 62844
Cp 1 2 3.009p
Rs 1 N3 0.298
L1 N3 2 48.357u
.ends 5848_784774156_56u
*******
.subckt 5848_784774168_68u 1 2
Rp 1 2 76697
Cp 1 2 3.081p
Rs 1 N3 0.313
L1 N3 2 59.979u
.ends 5848_784774168_68u
*******
.subckt 5848_784774182_82u 1 2
Rp 1 2 99452
Cp 1 2 3.405p
Rs 1 N3 0.475
L1 N3 2 74.566u
.ends 5848_784774182_82u
*******
.subckt 5848_78477420_100u 1 2
Rp 1 2 121927
Cp 1 2 3.348p
Rs 1 N3 0.51
L1 N3 2 90.852u
.ends 5848_78477420_100u
*******
.subckt 5848_784774212_120u 1 2
Rp 1 2 140140
Cp 1 2 3.348p
Rs 1 N3 0.66
L1 N3 2 102.363u
.ends 5848_784774212_120u
*******
.subckt 5848_784774215_150u 1 2
Rp 1 2 159467
Cp 1 2 3.482p
Rs 1 N3 0.72
L1 N3 2 130.131u
.ends 5848_784774215_150u
*******
.subckt 5848_784774218_180u 1 2
Rp 1 2 189610
Cp 1 2 3.247p
Rs 1 N3 0.85
L1 N3 2 167.071u
.ends 5848_784774218_180u
*******
.subckt 5848_784774222_220u 1 2
Rp 1 2 208937
Cp 1 2 3.388p
Rs 1 N3 0.945
L1 N3 2 195.681u
.ends 5848_784774222_220u
*******
.subckt 7850_784775022_2.2u 1 2
Rp 1 2 5325
Cp 1 2 2.151p
Rs 1 N3 0.008
L1 N3 2 1.889u
.ends 7850_784775022_2.2u
*******
.subckt 7850_784775047_4.7u 1 2
Rp 1 2 9103
Cp 1 2 2.498p
Rs 1 N3 0.016
L1 N3 2 3.751u
.ends 7850_784775047_4.7u
*******
.subckt 7850_784775056_5.6u 1 2
Rp 1 2 10274
Cp 1 2 2.738p
Rs 1 N3 0.018
L1 N3 2 4.375u
.ends 7850_784775056_5.6u
*******
.subckt 7850_784775068_6.8u 1 2
Rp 1 2 13545
Cp 1 2 2.723p
Rs 1 N3 0.022
L1 N3 2 5.769u
.ends 7850_784775068_6.8u
*******
.subckt 7850_784775082_8.2u 1 2
Rp 1 2 15056
Cp 1 2 3.046p
Rs 1 N3 0.024
L1 N3 2 6.629u
.ends 7850_784775082_8.2u
*******
.subckt 7850_78477510_10u 1 2
Rp 1 2 16424
Cp 1 2 2.779p
Rs 1 N3 0.04
L1 N3 2 8.061u
.ends 7850_78477510_10u
*******
.subckt 7850_784775112_12u 1 2
Rp 1 2 20036
Cp 1 2 3.195p
Rs 1 N3 0.042
L1 N3 2 9.631u
.ends 7850_784775112_12u
*******
.subckt 7850_784775115_15u 1 2
Rp 1 2 24297
Cp 1 2 3.216p
Rs 1 N3 0.044
L1 N3 2 13.006u
.ends 7850_784775115_15u
*******
.subckt 7850_784775118_18u 1 2
Rp 1 2 27614
Cp 1 2 3.321p
Rs 1 N3 0.053
L1 N3 2 15.149u
.ends 7850_784775118_18u
*******
.subckt 7850_784775122_22u 1 2
Rp 1 2 30904
Cp 1 2 3.29p
Rs 1 N3 0.065
L1 N3 2 17.549u
.ends 7850_784775122_22u
*******
.subckt 7850_784775127_27u 1 2
Rp 1 2 45613
Cp 1 2 3.55p
Rs 1 N3 0.074
L1 N3 2 22.657u
.ends 7850_784775127_27u
*******
.subckt 7850_784775133_33u 1 2
Rp 1 2 44853
Cp 1 2 3.438p
Rs 1 N3 0.089
L1 N3 2 28.459u
.ends 7850_784775133_33u
*******
.subckt 7850_784775139_39u 1 2
Rp 1 2 47106
Cp 1 2 3.639p
Rs 1 N3 0.116
L1 N3 2 31.967u
.ends 7850_784775139_39u
*******
.subckt 7850_784775147_47u 1 2
Rp 1 2 61345
Cp 1 2 13.35p
Rs 1 N3 0.134
L1 N3 2 33.411u
.ends 7850_784775147_47u
*******
.subckt 7850_784775168_68u 1 2
Rp 1 2 77918
Cp 1 2 3.664p
Rs 1 N3 0.218
L1 N3 2 58.886u
.ends 7850_784775168_68u
*******
.subckt 7850_784775182_82u 1 2
Rp 1 2 86377
Cp 1 2 3.867p
Rs 1 N3 0.248
L1 N3 2 71.757u
.ends 7850_784775182_82u
*******
.subckt 7850_78477520_100u 1 2
Rp 1 2 104821
Cp 1 2 3.713p
Rs 1 N3 0.281
L1 N3 2 82.03u
.ends 7850_78477520_100u
*******
.subckt 7850_784775212_120u 1 2
Rp 1 2 91873
Cp 1 2 20.977p
Rs 1 N3 0.34
L1 N3 2 99.003u
.ends 7850_784775212_120u
*******
.subckt 7850_784775215_150u 1 2
Rp 1 2 168654
Cp 1 2 3.941p
Rs 1 N3 0.467
L1 N3 2 128.415u
.ends 7850_784775215_150u
*******
.subckt 7850_784775218_180u 1 2
Rp 1 2 158858
Cp 1 2 4.027p
Rs 1 N3 0.574
L1 N3 2 168.879u
.ends 7850_784775218_180u
*******
.subckt 7850_784775222_220u 1 2
Rp 1 2 195165
Cp 1 2 3.728p
Rs 1 N3 0.614
L1 N3 2 194.368u
.ends 7850_784775222_220u
*******
.subckt 7850_784775227_270u 1 2
Rp 1 2 194699
Cp 1 2 4.392p
Rs 1 N3 0.699
L1 N3 2 224.595u
.ends 7850_784775227_270u
*******
.subckt 7850_784775233_330u 1 2
Rp 1 2 213144
Cp 1 2 4.501p
Rs 1 N3 0.98
L1 N3 2 260.153u
.ends 7850_784775233_330u
*******
.subckt 7850_784775239_390u 1 2
Rp 1 2 300959
Cp 1 2 3.983p
Rs 1 N3 1.151
L1 N3 2 364.959u
.ends 7850_784775239_390u
*******
.subckt 7850_784775247_470u 1 2
Rp 1 2 242537
Cp 1 2 4.045p
Rs 1 N3 1.37
L1 N3 2 400.519u
.ends 7850_784775247_470u
*******
