**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  Aluminum Electrolytic Capacitors
* Matchcode:              WCAP-AS5H
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/20/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 865230640004_470nF 1 2
Rser 1 3 2.47418974398
Lser 2 4 1.492372247E-09
C1 3 4 0.00000047
Rpar 3 4 16666666.6666667
.ends 865230640004_470nF
*******
.subckt 865230640005_1uF 1 2
Rser 1 3 2.66794645225
Lser 2 4 8.51832959E-10
C1 3 4 0.000001
Rpar 3 4 16666666.6666667
.ends 865230640005_1uF
*******
.subckt 865230640006_2.2uF 1 2
Rser 1 3 2.2608421566
Lser 2 4 1.3849563E-09
C1 3 4 0.0000022
Rpar 3 4 16666666.6666667
.ends 865230640006_2.2uF
*******
.subckt 865230640007_3.3uF 1 2
Rser 1 3 2.68570511593
Lser 2 4 9.96555496E-10
C1 3 4 0.0000033
Rpar 3 4 16666666.6666667
.ends 865230640007_3.3uF
*******
.subckt 865230440001_4.7uF 1 2
Rser 1 3 1.5
Lser 2 4 0.00000000000055
C1 3 4 0.0000047
Rpar 3 4 8333333.33333333
.ends 865230440001_4.7uF
*******
.subckt 865230540001_4.7uF 1 2
Rser 1 3 2.49723366161
Lser 2 4 1.483332833E-09
C1 3 4 0.0000047
Rpar 3 4 11666666.6666667
.ends 865230540001_4.7uF
*******
.subckt 865230340001_10uF 1 2
Rser 1 3 2.29118477444
Lser 2 4 1.062989445E-09
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 865230340001_10uF
*******
.subckt 865230440002_10uF 1 2
Rser 1 3 1.95
Lser 2 4 0.00000000000007
C1 3 4 0.00001
Rpar 3 4 8333333.33333333
.ends 865230440002_10uF
*******
.subckt 865230140001_22uF 1 2
Rser 1 3 2.4262199213
Lser 2 4 9.63393805E-10
C1 3 4 0.000022
Rpar 3 4 2100000
.ends 865230140001_22uF
*******
.subckt 865230642008_4.7uF 1 2
Rser 1 3 1.74334241586
Lser 2 4 2.808642261E-09
C1 3 4 0.0000047
Rpar 3 4 16666666.6666667
.ends 865230642008_4.7uF
*******
.subckt 865230542002_10uF 1 2
Rser 1 3 1.62310107626
Lser 2 4 2.55094298E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865230542002_10uF
*******
.subckt 865230342002_22uF 1 2
Rser 1 3 1.63827766347
Lser 2 4 1.77818178E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865230342002_22uF
*******
.subckt 865230242001_22uF 1 2
Rser 1 3 1.59163089519
Lser 2 4 2.782802747E-09
C1 3 4 0.000022
Rpar 3 4 3333333.33333333
.ends 865230242001_22uF
*******
.subckt 865230142002_33uF 1 2
Rser 1 3 1.46979022371
Lser 2 4 2.843754388E-09
C1 3 4 0.000033
Rpar 3 4 2100000
.ends 865230142002_33uF
*******
.subckt 865230242002_33uF 1 2
Rser 1 3 1.61907751429
Lser 2 4 0.000000001824
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865230242002_33uF
*******
.subckt 865230142003_47uF 1 2
Rser 1 3 1.35945323523
Lser 2 4 2.492556603E-09
C1 3 4 0.000047
Rpar 3 4 2100000
.ends 865230142003_47uF
*******
.subckt 865230643009_10uF 1 2
Rser 1 3 1.15848603831
Lser 2 4 2.253179561E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865230643009_10uF
*******
.subckt 865230443003_22uF 1 2
Rser 1 3 0.61
Lser 2 4 0.0000000001
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865230443003_22uF
*******
.subckt 865230645010_22uF 1 2
Rser 1 3 0.64433896064
Lser 2 4 4.11393679E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865230645010_22uF
*******
.subckt 865230543003_22uF 1 2
Rser 1 3 0.75722878803
Lser 2 4 3.831409158E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 865230543003_22uF
*******
.subckt 865230343003_33uF 1 2
Rser 1 3 0.794148504904
Lser 2 4 4.036746464E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865230343003_33uF
*******
.subckt 865230545004_33uF 1 2
Rser 1 3 0.647354185398
Lser 2 4 4.427850728E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865230545004_33uF
*******
.subckt 865230443004_33uF 1 2
Rser 1 3 0.61
Lser 2 4 0.000000000076
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865230443004_33uF
*******
.subckt 865230343004_47uF 1 2
Rser 1 3 0.801370085672
Lser 2 4 4.120619727E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865230343004_47uF
*******
.subckt 865230445005_47uF 1 2
Rser 1 3 0.38
Lser 2 4 0.0000000002
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865230445005_47uF
*******
.subckt 865230243003_47uF 1 2
Rser 1 3 0.811054859702
Lser 2 4 4.070325673E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865230243003_47uF
*******
.subckt 865230345005_100uF 1 2
Rser 1 3 0.488
Lser 2 4 2.808093044E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865230345005_100uF
*******
.subckt 865230143004_100uF 1 2
Rser 1 3 0.8503949862
Lser 2 4 3.796940524E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865230143004_100uF
*******
.subckt 865230245004_100uF 1 2
Rser 1 3 0.327
Lser 2 4 2.719633456E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865230245004_100uF
*******
.subckt 865230145005_220uF 1 2
Rser 1 3 0.285
Lser 2 4 0.00000000013
C1 3 4 0.00022
Rpar 3 4 454545.454545454
.ends 865230145005_220uF
*******
.subckt 865230364011_220uF 1 2
Rser 1 3 0.28
Lser 2 4 0.00000000235
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865230364011_220uF
*******
.subckt 865230653011_33uF 1 2
Rser 1 3 0.575738257859
Lser 2 4 4.960298117E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865230653011_33uF
*******
.subckt 865230653012_47uF 1 2
Rser 1 3 0.336814650022
Lser 2 4 5.079815563E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865230653012_47uF
*******
.subckt 865230553005_47uF 1 2
Rser 1 3 0.35687838853
Lser 2 4 5.202348961E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865230553005_47uF
*******
.subckt 865230453006_100uF 1 2
Rser 1 3 0.169
Lser 2 4 5.16204113085425E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865230453006_100uF
*******
.subckt 865230253005_220uF 1 2
Rser 1 3 0.215
Lser 2 4 0.0000000004
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865230253005_220uF
*******
.subckt 865230153006_330uF 1 2
Rser 1 3 0.22518
Lser 2 4 3.886945652E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865230153006_330uF
*******
.subckt 865230657013_100uF 1 2
Rser 1 3 0.189
Lser 2 4 5.72884434804354E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865230657013_100uF
*******
.subckt 865230557006_100uF 1 2
Rser 1 3 0.135
Lser 2 4 0.0000000015
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865230557006_100uF
*******
.subckt 865230357006_220uF 1 2
Rser 1 3 0.15
Lser 2 4 0.0000000013
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865230357006_220uF
*******
.subckt 865230457007_220uF 1 2
Rser 1 3 0.107
Lser 2 4 0.0000000011
C1 3 4 0.00022
Rpar 3 4 454545.454545454
.ends 865230457007_220uF
*******
.subckt 865230557007_220uF 1 2
Rser 1 3 0.115
Lser 2 4 0.0000000013
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865230557007_220uF
*******
.subckt 865230357007_330uF 1 2
Rser 1 3 0.097
Lser 2 4 6.82551885070387E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865230357007_330uF
*******
.subckt 865230457008_330uF 1 2
Rser 1 3 0.08
Lser 2 4 0.0000000014
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865230457008_330uF
*******
.subckt 865230257006_330uF 1 2
Rser 1 3 0.095
Lser 2 4 0.000000001
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865230257006_330uF
*******
.subckt 865230657014_330uF 1 2
Rser 1 3 0.085
Lser 2 4 0.0000000013
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865230657014_330uF
*******
.subckt 865230357008_470uF 1 2
Rser 1 3 0.087
Lser 2 4 0.0000000008
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865230357008_470uF
*******
.subckt 865230157007_470uF 1 2
Rser 1 3 0.1
Lser 2 4 0.0000000007
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865230157007_470uF
*******
.subckt 865230257007_470uF 1 2
Rser 1 3 0.09
Lser 2 4 0.000000001
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865230257007_470uF
*******
.subckt 865230157008_1mF 1 2
Rser 1 3 0.107
Lser 2 4 0.0000000007
C1 3 4 0.001
Rpar 3 4 100000
.ends 865230157008_1mF
*******
