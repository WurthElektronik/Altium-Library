**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  MLCCs - Multilayer Ceramic Chip Capacitors
* Matchcode:              WCAP-CSGP_10V
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/20/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0201_885012204005_10nF 1 2
Rser 1 3 0.0631
Lser 2 4 0.000000000217
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012204005_10nF
*******
.subckt 0201_885012104012_10nF 1 2
Rser 1 3 0.0632
Lser 2 4 0.000000000213
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012104012_10nF
*******
.subckt 0201_885012104013_47nF 1 2
Rser 1 3 0.06035
Lser 2 4 0.00000000022
C1 3 4 0.000000047
Rpar 3 4 2000000000
.ends 0201_885012104013_47nF
*******
.subckt 0201_885012104002_100nF 1 2
Rser 1 3 0.02596
Lser 2 4 0.00000000018
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0201_885012104002_100nF
*******
.subckt 0201_885012104006_220nF 1 2
Rser 1 3 0.02291
Lser 2 4 0.00000000015
C1 3 4 0.00000022
Rpar 3 4 200000000
.ends 0201_885012104006_220nF
*******
.subckt 0402_885012005001_1pF 1 2
Rser 1 3 1.871
Lser 2 4 0.00000000033
C1 3 4 0.000000000001
Rpar 3 4 10000000000
.ends 0402_885012005001_1pF
*******
.subckt 0402_885012005002_1.5pF 1 2
Rser 1 3 0.9
Lser 2 4 0.00000000031
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0402_885012005002_1.5pF
*******
.subckt 0402_885012005004_3.3pF 1 2
Rser 1 3 0.7
Lser 2 4 0.00000000039
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0402_885012005004_3.3pF
*******
.subckt 0402_885012005005_4.7pF 1 2
Rser 1 3 1
Lser 2 4 0.00000000041
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0402_885012005005_4.7pF
*******
.subckt 0402_885012005006_6.8pF 1 2
Rser 1 3 0.4886
Lser 2 4 0.00000000032
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0402_885012005006_6.8pF
*******
.subckt 0402_885012005007_10pF 1 2
Rser 1 3 0.494547705824
Lser 2 4 3.67389142E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005007_10pF
*******
.subckt 0402_885012005008_15pF 1 2
Rser 1 3 0.388190780491
Lser 2 4 3.17307789E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885012005008_15pF
*******
.subckt 0402_885012005009_22pF 1 2
Rser 1 3 0.316230222598
Lser 2 4 2.88077478E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885012005009_22pF
*******
.subckt 0402_885012005010_33pF 1 2
Rser 1 3 0.249324470259
Lser 2 4 2.84730223E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005010_33pF
*******
.subckt 0402_885012005011_47pF 1 2
Rser 1 3 0.235686289563
Lser 2 4 2.78272514E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005011_47pF
*******
.subckt 0402_885012005012_68pF 1 2
Rser 1 3 0.188011183755
Lser 2 4 2.62979806E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005012_68pF
*******
.subckt 0402_885012005013_100pF 1 2
Rser 1 3 0.145490051878
Lser 2 4 2.5124412E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005013_100pF
*******
.subckt 0402_885012005014_150pF 1 2
Rser 1 3 0.102893245885
Lser 2 4 2.1894381E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012005014_150pF
*******
.subckt 0402_885012005015_220pF 1 2
Rser 1 3 0.0932691679838
Lser 2 4 1.50271806E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012005015_220pF
*******
.subckt 0402_885012005016_330pF 1 2
Rser 1 3 0.0893241489871
Lser 2 4 3.29295953E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012005016_330pF
*******
.subckt 0402_885012005017_470pF 1 2
Rser 1 3 0.0149178531097
Lser 2 4 3.26241368E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012005017_470pF
*******
.subckt 0402_885012005018_1nF 1 2
Rser 1 3 0.0157004412396
Lser 2 4 3.37941862E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012005018_1nF
*******
.subckt 0402_885012105009_68nF 1 2
Rser 1 3 0.0638704519417
Lser 2 4 2.20630867E-10
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0402_885012105009_68nF
*******
.subckt 0402_885012105010_100nF 1 2
Rser 1 3 0.0268043216773
Lser 2 4 3.11178988E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012105010_100nF
*******
.subckt 0402_885012105011_220nF 1 2
Rser 1 3 0.0122717751401
Lser 2 4 3.48439745E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0402_885012105011_220nF
*******
.subckt 0402_885012105012_1uF 1 2
Rser 1 3 0.00986403339919
Lser 2 4 3.2821055E-10
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0402_885012105012_1uF
*******
.subckt 0402_885012105013_2.2uF 1 2
Rser 1 3 0.019
Lser 2 4 0.000000001
C1 3 4 0.0000022
Rpar 3 4 20000000
.ends 0402_885012105013_2.2uF
*******
.subckt 0402_885012205001_100pF 1 2
Rser 1 3 0.78619
Lser 2 4 0.00000000015138
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012205001_100pF
*******
.subckt 0402_885012205002_220pF 1 2
Rser 1 3 0.5727
Lser 2 4 1.77695991E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012205002_220pF
*******
.subckt 0402_885012205003_330pF 1 2
Rser 1 3 0.43753
Lser 2 4 0.00000000020201
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012205003_330pF
*******
.subckt 0402_885012205004_470pF 1 2
Rser 1 3 0.33537
Lser 2 4 0.00000000018013
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012205004_470pF
*******
.subckt 0402_885012205005_680pF 1 2
Rser 1 3 0.26133
Lser 2 4 0.00000000015756
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0402_885012205005_680pF
*******
.subckt 0402_885012205006_1nF 1 2
Rser 1 3 0.19089
Lser 2 4 0.00000000017743
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205006_1nF
*******
.subckt 0402_885012205007_1.5nF 1 2
Rser 1 3 0.16721
Lser 2 4 0.00000000024076
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0402_885012205007_1.5nF
*******
.subckt 0402_885012205008_2.2nF 1 2
Rser 1 3 0.11524
Lser 2 4 0.000000000227222
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0402_885012205008_2.2nF
*******
.subckt 0402_885012205009_3.3nF 1 2
Rser 1 3 0.0897
Lser 2 4 0.00000000023518
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0402_885012205009_3.3nF
*******
.subckt 0402_885012205010_4.7nF 1 2
Rser 1 3 0.05632
Lser 2 4 0.00000000018931
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205010_4.7nF
*******
.subckt 0402_885012205011_6.8nF 1 2
Rser 1 3 0.04164
Lser 2 4 0.00000000021064
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0402_885012205011_6.8nF
*******
.subckt 0402_885012205012_10nF 1 2
Rser 1 3 0.0531398956639
Lser 2 4 0.00000000022
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0402_885012205012_10nF
*******
.subckt 0402_885012205013_15nF 1 2
Rser 1 3 0.03039
Lser 2 4 0.00000000022583
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0402_885012205013_15nF
*******
.subckt 0402_885012205014_22nF 1 2
Rser 1 3 0.01645
Lser 2 4 0.00000000020049
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0402_885012205014_22nF
*******
.subckt 0402_885012205015_33nF 1 2
Rser 1 3 0.00701
Lser 2 4 0.00000000023581
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0402_885012205015_33nF
*******
.subckt 0402_885012205016_47nF 1 2
Rser 1 3 0.0071
Lser 2 4 0.0000000002065
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0402_885012205016_47nF
*******
.subckt 0402_885012205017_68nF 1 2
Rser 1 3 0.01539
Lser 2 4 0.00000000023044
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0402_885012205017_68nF
*******
.subckt 0402_885012205018_100nF 1 2
Rser 1 3 0.0183525691398
Lser 2 4 3.07541467E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205018_100nF
*******
.subckt 0402_885012105026_4.7uF 1 2
Rser 1 3 0.00852
Lser 2 4 0.000000001132
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0402_885012105026_4.7uF
*******
.subckt 0603_885012006001_4.7pF 1 2
Rser 1 3 0.307143942354
Lser 2 4 3.18870536E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0603_885012006001_4.7pF
*******
.subckt 0603_885012006002_10pF 1 2
Rser 1 3 0.668
Lser 2 4 0.00000000056
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006002_10pF
*******
.subckt 0603_885012006003_15pF 1 2
Rser 1 3 0.318625808147
Lser 2 4 7.07424269E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006003_15pF
*******
.subckt 0603_885012006004_22pF 1 2
Rser 1 3 0.34819611654
Lser 2 4 7.75018519E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006004_22pF
*******
.subckt 0603_885012006005_33pF 1 2
Rser 1 3 0.266845513997
Lser 2 4 8.03723788E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006005_33pF
*******
.subckt 0603_885012006006_47pF 1 2
Rser 1 3 0.196782783005
Lser 2 4 7.59426691E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006006_47pF
*******
.subckt 0603_885012006007_68pF 1 2
Rser 1 3 0.153641735222
Lser 2 4 7.22489136E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006007_68pF
*******
.subckt 0603_885012006008_100pF 1 2
Rser 1 3 0.110129832129
Lser 2 4 6.73785263E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006008_100pF
*******
.subckt 0603_885012006009_150pF 1 2
Rser 1 3 0.0793891689318
Lser 2 4 6.22415559E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006009_150pF
*******
.subckt 0603_885012006010_220pF 1 2
Rser 1 3 0.088220302088
Lser 2 4 6.95492511E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012006010_220pF
*******
.subckt 0603_885012006011_330pF 1 2
Rser 1 3 0.0993151086205
Lser 2 4 4.18653134E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006011_330pF
*******
.subckt 0603_885012006012_470pF 1 2
Rser 1 3 0.0757443435992
Lser 2 4 3.66481782E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006012_470pF
*******
.subckt 0603_885012006013_680pF 1 2
Rser 1 3 0.0602766942369
Lser 2 4 3.26882078E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006013_680pF
*******
.subckt 0603_885012006014_1nF 1 2
Rser 1 3 0.0434067925003
Lser 2 4 4.09321859E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006014_1nF
*******
.subckt 0603_885012006015_2.2nF 1 2
Rser 1 3 0.0307077888885
Lser 2 4 3.39702907E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012006015_2.2nF
*******
.subckt 0603_885012006016_3.3nF 1 2
Rser 1 3 0.0275317919224
Lser 2 4 3.37901927E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012006016_3.3nF
*******
.subckt 0603_885012106007_330nF 1 2
Rser 1 3 0.0111038975002
Lser 2 4 3.20933284E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012106007_330nF
*******
.subckt 0603_885012106008_470nF 1 2
Rser 1 3 0.00949633292517
Lser 2 4 2.70539302E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0603_885012106008_470nF
*******
.subckt 0603_885012106009_680nF 1 2
Rser 1 3 0.0112015362567
Lser 2 4 3.50610132E-10
C1 3 4 0.00000068
Rpar 3 4 200000000
.ends 0603_885012106009_680nF
*******
.subckt 0603_885012106010_1uF 1 2
Rser 1 3 0.00802031801588
Lser 2 4 3.00240209E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012106010_1uF
*******
.subckt 0603_885012106011_2.2uF 1 2
Rser 1 3 0.00618507884481
Lser 2 4 2.53136283E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0603_885012106011_2.2uF
*******
.subckt 0603_885012106012_4.7uF 1 2
Rser 1 3 0.00455496693599
Lser 2 4 5.03384516E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0603_885012106012_4.7uF
*******
.subckt 0603_885012206003_100pF 1 2
Rser 1 3 0.86219
Lser 2 4 0.00000000020992
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206003_100pF
*******
.subckt 0603_885012206004_220pF 1 2
Rser 1 3 0.55667
Lser 2 4 0.00000000030069
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012206004_220pF
*******
.subckt 0603_885012206005_330pF 1 2
Rser 1 3 0.43756
Lser 2 4 0.00000000026062
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206005_330pF
*******
.subckt 0603_885012206006_470pF 1 2
Rser 1 3 0.37246
Lser 2 4 0.00000000030107
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206006_470pF
*******
.subckt 0603_885012206007_680pF 1 2
Rser 1 3 0.31851
Lser 2 4 0.00000000040239
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206007_680pF
*******
.subckt 0603_885012206008_1nF 1 2
Rser 1 3 0.24958
Lser 2 4 0.00000000040399
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206008_1nF
*******
.subckt 0603_885012206009_1.5nF 1 2
Rser 1 3 0.20086
Lser 2 4 0.00000000033824
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206009_1.5nF
*******
.subckt 0603_885012206010_2.2nF 1 2
Rser 1 3 0.14948
Lser 2 4 0.00000000033334
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012206010_2.2nF
*******
.subckt 0603_885012206011_3.3nF 1 2
Rser 1 3 0.12415
Lser 2 4 0.00000000032537
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206011_3.3nF
*******
.subckt 0603_885012206012_4.7nF 1 2
Rser 1 3 0.07518
Lser 2 4 0.0000000003009
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206012_4.7nF
*******
.subckt 0603_885012206013_6.8nF 1 2
Rser 1 3 0.07031
Lser 2 4 0.00000000039053
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206013_6.8nF
*******
.subckt 0603_885012206014_10nF 1 2
Rser 1 3 0.04641
Lser 2 4 0.00000000025735
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206014_10nF
*******
.subckt 0603_885012206015_15nF 1 2
Rser 1 3 0.03908
Lser 2 4 0.00000000026071
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0603_885012206015_15nF
*******
.subckt 0603_885012206016_22nF 1 2
Rser 1 3 0.02302
Lser 2 4 0.00000000023719
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885012206016_22nF
*******
.subckt 0603_885012206017_33nF 1 2
Rser 1 3 0.01243
Lser 2 4 0.00000000025982
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0603_885012206017_33nF
*******
.subckt 0603_885012206018_47nF 1 2
Rser 1 3 0.01343
Lser 2 4 0.00000000024476
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0603_885012206018_47nF
*******
.subckt 0603_885012206019_68nF 1 2
Rser 1 3 0.0155
Lser 2 4 0.00000000030737
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0603_885012206019_68nF
*******
.subckt 0603_885012206020_100nF 1 2
Rser 1 3 0.0188883213835
Lser 2 4 4.53593763E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206020_100nF
*******
.subckt 0603_885012206021_150nF 1 2
Rser 1 3 0.0221138242279
Lser 2 4 4.07625742E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0603_885012206021_150nF
*******
.subckt 0603_885012206022_220nF 1 2
Rser 1 3 0.0146862228843
Lser 2 4 4.43010481E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012206022_220nF
*******
.subckt 0603_885012206023_330nF 1 2
Rser 1 3 0.0113479919005
Lser 2 4 4.48567636E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012206023_330nF
*******
.subckt 0603_885012206024_470nF 1 2
Rser 1 3 0.00961049589993
Lser 2 4 4.09343651E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0603_885012206024_470nF
*******
.subckt 0603_885012206025_680nF 1 2
Rser 1 3 0.00730055384166
Lser 2 4 4.35162169E-10
C1 3 4 0.00000068
Rpar 3 4 200000000
.ends 0603_885012206025_680nF
*******
.subckt 0603_885012206026_1uF 1 2
Rser 1 3 0.00743560640346
Lser 2 4 2.29632839E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012206026_1uF
*******
.subckt 0603_885012206027_2.2uF 1 2
Rser 1 3 0.00844425861819
Lser 2 4 2.90335669E-10
C1 3 4 0.0000022
Rpar 3 4 20000000
.ends 0603_885012206027_2.2uF
*******
.subckt 0603_885012106032_22uF 1 2
Rser 1 3 0.0055
Lser 2 4 0.0000000008
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 0603_885012106032_22uF
*******
.subckt 0805_885012007001_15pF 1 2
Rser 1 3 0.322686614764
Lser 2 4 5.17792028E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007001_15pF
*******
.subckt 0805_885012007002_22pF 1 2
Rser 1 3 0.304017782882
Lser 2 4 6.06807592E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0805_885012007002_22pF
*******
.subckt 0805_885012007003_33pF 1 2
Rser 1 3 0.278413141435
Lser 2 4 5.73322702E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007003_33pF
*******
.subckt 0805_885012007004_100pF 1 2
Rser 1 3 0.144376756
Lser 2 4 4.19735168E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007004_100pF
*******
.subckt 0805_885012007005_150pF 1 2
Rser 1 3 0.132070069125
Lser 2 4 4.14007712E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007005_150pF
*******
.subckt 0805_885012007006_330pF 1 2
Rser 1 3 0.0858219234392
Lser 2 4 4.4258651E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007006_330pF
*******
.subckt 0805_885012007007_470pF 1 2
Rser 1 3 0.0754569114616
Lser 2 4 4.35286885E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007007_470pF
*******
.subckt 0805_885012007008_1nF 1 2
Rser 1 3 0.0525130505561
Lser 2 4 4.16381481E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007008_1nF
*******
.subckt 0805_885012007009_10nF 1 2
Rser 1 3 0.0143302506767
Lser 2 4 2.53788056E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012007009_10nF
*******
.subckt 0805_885012107007_2.2uF 1 2
Rser 1 3 0.00451361812717
Lser 2 4 2.56807852E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012107007_2.2uF
*******
.subckt 0805_885012107008_3.3uF 1 2
Rser 1 3 0.00416445411098
Lser 2 4 3.00167169E-10
C1 3 4 0.0000033
Rpar 3 4 30000000
.ends 0805_885012107008_3.3uF
*******
.subckt 0805_885012107009_4.7uF 1 2
Rser 1 3 0.00333037459922
Lser 2 4 2.41667028E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0805_885012107009_4.7uF
*******
.subckt 0805_885012107010_10uF 1 2
Rser 1 3 0.00257315295813
Lser 2 4 4.16651033E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 0805_885012107010_10uF
*******
.subckt 0805_885012107011_22uF 1 2
Rser 1 3 0.00309713657007
Lser 2 4 2.86347556E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 0805_885012107011_22uF
*******
.subckt 0805_885012207004_100pF 1 2
Rser 1 3 0.88264
Lser 2 4 0.00000000031858
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207004_100pF
*******
.subckt 0805_885012207005_220pF 1 2
Rser 1 3 0.50995
Lser 2 4 0.00000000027274
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012207005_220pF
*******
.subckt 0805_885012207006_470pF 1 2
Rser 1 3 0.31274
Lser 2 4 0.00000000031898
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207006_470pF
*******
.subckt 0805_885012207007_1nF 1 2
Rser 1 3 0.1905
Lser 2 4 0.00000000028002
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207007_1nF
*******
.subckt 0805_885012207008_1.5nF 1 2
Rser 1 3 0.16519
Lser 2 4 0.00000000038865
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207008_1.5nF
*******
.subckt 0805_885012207009_2.2nF 1 2
Rser 1 3 0.02478
Lser 2 4 0.00000000027522
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012207009_2.2nF
*******
.subckt 0805_885012207010_3.3nF 1 2
Rser 1 3 0.02239
Lser 2 4 0.00000000023565
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207010_3.3nF
*******
.subckt 0805_885012207011_10nF 1 2
Rser 1 3 0.04883
Lser 2 4 0.00000000031494
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207011_10nF
*******
.subckt 0805_885012207012_15nF 1 2
Rser 1 3 0.0512
Lser 2 4 0.00000000030048
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0805_885012207012_15nF
*******
.subckt 0805_885012207013_22nF 1 2
Rser 1 3 0.03858
Lser 2 4 0.00000000031876
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0805_885012207013_22nF
*******
.subckt 0805_885012207014_33nF 1 2
Rser 1 3 0.03079
Lser 2 4 0.00000000030588
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0805_885012207014_33nF
*******
.subckt 0805_885012207015_47nF 1 2
Rser 1 3 0.02162
Lser 2 4 0.0000000002672
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0805_885012207015_47nF
*******
.subckt 0805_885012207016_100nF 1 2
Rser 1 3 0.0162501221785
Lser 2 4 0.000000000375
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207016_100nF
*******
.subckt 0805_885012207017_150nF 1 2
Rser 1 3 0.0143154309487
Lser 2 4 4.47033542E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0805_885012207017_150nF
*******
.subckt 0805_885012207018_220nF 1 2
Rser 1 3 0.0114343175461
Lser 2 4 4.37838091E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885012207018_220nF
*******
.subckt 0805_885012207019_330nF 1 2
Rser 1 3 0.0106449562538
Lser 2 4 4.87419012E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885012207019_330nF
*******
.subckt 0805_885012207020_470nF 1 2
Rser 1 3 0.00823353483639
Lser 2 4 4.7697612E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0805_885012207020_470nF
*******
.subckt 0805_885012207021_680nF 1 2
Rser 1 3 0.00756100048721
Lser 2 4 5.19694932E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0805_885012207021_680nF
*******
.subckt 0805_885012207022_1uF 1 2
Rser 1 3 0.00779960743902
Lser 2 4 2.50116995E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885012207022_1uF
*******
.subckt 0805_885012207023_1.5uF 1 2
Rser 1 3 0.00625640838813
Lser 2 4 3.16162321E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 0805_885012207023_1.5uF
*******
.subckt 0805_885012207024_2.2uF 1 2
Rser 1 3 0.00498465718149
Lser 2 4 2.58299749E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012207024_2.2uF
*******
.subckt 0805_885012207025_4.7uF 1 2
Rser 1 3 0.008
Lser 2 4 0.0000000006
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0805_885012207025_4.7uF
*******
.subckt 0805_885012207026_10uF 1 2
Rser 1 3 0.00369416302331
Lser 2 4 5.01488494E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0805_885012207026_10uF
*******
.subckt 1206_885012008001_10pF 1 2
Rser 1 3 0.446014275484
Lser 2 4 5.73571915E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1206_885012008001_10pF
*******
.subckt 1206_885012008002_22pF 1 2
Rser 1 3 0.299003095867
Lser 2 4 5.45254376E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1206_885012008002_22pF
*******
.subckt 1206_885012008003_47pF 1 2
Rser 1 3 0.21040740508
Lser 2 4 5.6609278E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885012008003_47pF
*******
.subckt 1206_885012008004_100pF 1 2
Rser 1 3 0.167865253643
Lser 2 4 4.85486348E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008004_100pF
*******
.subckt 1206_885012008005_470pF 1 2
Rser 1 3 0.115247377385
Lser 2 4 4.7229295E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012008005_470pF
*******
.subckt 1206_885012008006_2.2nF 1 2
Rser 1 3 0.0350339469969
Lser 2 4 1.042313537E-09
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012008006_2.2nF
*******
.subckt 1206_885012008007_6.8nF 1 2
Rser 1 3 0.0298615638448
Lser 2 4 9.14635803E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008007_6.8nF
*******
.subckt 1206_885012008008_10nF 1 2
Rser 1 3 0.0249778783357
Lser 2 4 9.13131263E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008008_10nF
*******
.subckt 1206_885012008009_22nF 1 2
Rser 1 3 0.011442234975
Lser 2 4 8.6240711E-10
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1206_885012008009_22nF
*******
.subckt 1206_885012008010_33nF 1 2
Rser 1 3 0.0092860021616
Lser 2 4 8.63894198E-10
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1206_885012008010_33nF
*******
.subckt 1206_885012108006_2.2uF 1 2
Rser 1 3 0.00715208568262
Lser 2 4 5.64041345E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012108006_2.2uF
*******
.subckt 1206_885012108007_3.3uF 1 2
Rser 1 3 0.00529476260464
Lser 2 4 6.12367847E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012108007_3.3uF
*******
.subckt 1206_885012108008_4.7uF 1 2
Rser 1 3 0.00610205096672
Lser 2 4 5.17669274E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012108008_4.7uF
*******
.subckt 1206_885012108009_6.8uF 1 2
Rser 1 3 0.00416216687199
Lser 2 4 6.95534046E-10
C1 3 4 0.0000068
Rpar 3 4 20000000
.ends 1206_885012108009_6.8uF
*******
.subckt 1206_885012108010_10uF 1 2
Rser 1 3 0.00362327531378
Lser 2 4 0.0000000008
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1206_885012108010_10uF
*******
.subckt 1206_885012108011_22uF 1 2
Rser 1 3 0.00240452659004
Lser 2 4 8.37875791E-10
C1 3 4 0.000022
Rpar 3 4 5000000
.ends 1206_885012108011_22uF
*******
.subckt 1206_885012108012_47uF 1 2
Rser 1 3 0.0027428064885
Lser 2 4 0.0000000008
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1206_885012108012_47uF
*******
.subckt 1206_885012208004_330pF 1 2
Rser 1 3 0.46442
Lser 2 4 0.00000000041059
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012208004_330pF
*******
.subckt 1206_885012208005_470pF 1 2
Rser 1 3 0.38435
Lser 2 4 0.00000000043066
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208005_470pF
*******
.subckt 1206_885012208006_1nF 1 2
Rser 1 3 0.22561
Lser 2 4 0.00000000045042
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208006_1nF
*******
.subckt 1206_885012208007_4.7nF 1 2
Rser 1 3 0.13666
Lser 2 4 0.00000000045064
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208007_4.7nF
*******
.subckt 1206_885012208008_10nF 1 2
Rser 1 3 0.06965
Lser 2 4 0.00000000068939
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208008_10nF
*******
.subckt 1206_885012208009_100nF 1 2
Rser 1 3 0.0244803326156
Lser 2 4 6.58788173E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885012208009_100nF
*******
.subckt 1206_885012208010_330nF 1 2
Rser 1 3 0.0123317635994
Lser 2 4 6.03276395E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1206_885012208010_330nF
*******
.subckt 1206_885012208011_470nF 1 2
Rser 1 3 0.010415539685
Lser 2 4 7.51451536E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1206_885012208011_470nF
*******
.subckt 1206_885012208012_680nF 1 2
Rser 1 3 0.00703741199294
Lser 2 4 7.17949052E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1206_885012208012_680nF
*******
.subckt 1206_885012208013_1uF 1 2
Rser 1 3 0.00648320483926
Lser 2 4 5.4243262E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885012208013_1uF
*******
.subckt 1206_885012208014_1.5uF 1 2
Rser 1 3 0.00911925278109
Lser 2 4 6.57782928E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 1206_885012208014_1.5uF
*******
.subckt 1206_885012208015_2.2uF 1 2
Rser 1 3 0.00662951285801
Lser 2 4 5.30235159E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012208015_2.2uF
*******
.subckt 1206_885012208016_3.3uF 1 2
Rser 1 3 0.00509978680029
Lser 2 4 6.27645723E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012208016_3.3uF
*******
.subckt 1206_885012208017_4.7uF 1 2
Rser 1 3 0.00357416297194
Lser 2 4 4.72459357E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012208017_4.7uF
*******
.subckt 1206_885012208018_10uF 1 2
Rser 1 3 0.00288901435933
Lser 2 4 7.48356777E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1206_885012208018_10uF
*******
.subckt 1206_885012208019_22uF 1 2
Rser 1 3 0.00343100506851
Lser 2 4 5.00393923E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1206_885012208019_22uF
*******
.subckt 1210_885012109005_10uF 1 2
Rser 1 3 0.00250479636867
Lser 2 4 7.49918881E-10
C1 3 4 0.00001
Rpar 3 4 50000000
.ends 1210_885012109005_10uF
*******
.subckt 1210_885012109006_22uF 1 2
Rser 1 3 0.00272955719838
Lser 2 4 9.31961125E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1210_885012109006_22uF
*******
.subckt 1210_885012109007_47uF 1 2
Rser 1 3 0.00210105515092
Lser 2 4 0.0000000009
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1210_885012109007_47uF
*******
.subckt 1210_885012209001_47nF 1 2
Rser 1 3 0.03203
Lser 2 4 0.00000000012248
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1210_885012209001_47nF
*******
.subckt 1210_885012209002_220nF 1 2
Rser 1 3 0.0108946736088
Lser 2 4 5.13453415E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1210_885012209002_220nF
*******
.subckt 1210_885012209003_1uF 1 2
Rser 1 3 0.00441457708348
Lser 2 4 3.73414796E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209003_1uF
*******
.subckt 1210_885012209004_4.7uF 1 2
Rser 1 3 0.0051217091228
Lser 2 4 5.20978006E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012209004_4.7uF
*******
.subckt 1210_885012209005_10uF 1 2
Rser 1 3 0.00237372157538
Lser 2 4 7.95583466E-10
C1 3 4 0.00001
Rpar 3 4 100000000
.ends 1210_885012209005_10uF
*******
.subckt 1210_885012209006_22uF 1 2
Rser 1 3 0.0039
Lser 2 4 0.00000000075
C1 3 4 0.000022
Rpar 3 4 10000000
.ends 1210_885012209006_22uF
*******
