**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Common Mode Power Line Choke Nanocrystalline 
* Matchcode:              WE-CMBNC 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-26
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.SUBCKT CMBNC  1  2  3  4  PARAMS:
+  L1=0.00060538
+  L2=0.00010035
+  L3=0.00004247
+  L4=0.00001022
+  L5=0.000000036
+  C1=0.000000000003
+  C2=0.000000000001
+  RS1=8828
+  RS2=1447
+  RS3=703
+  RS4=678
+  RS5=509
+  R2=0.11
+  DL3=0.00000031037
+  DL4=0.00000001106
+  DC3=0.00000000000019056
+  DC4=0.000000000007
+  DR3=1000
+  DR4=4500
+  DR5=11000
+  DR6=438
+  Rdc=0.43
+  ck=12.5pF
L5  N010  N009  {L3}
R50  N010  N009  {Rs3}
C3  N500  N001  {C1}
R500  4  N500  {R2}
L1  4  N011  {L1}
R51  4  N011  {Rs1}
L3  N011  N010  {L2}
R52  N011  N010  {Rs2}
L6  N014  N013  {L3}
R53  N014  N013  {Rs3}
C4  N501  N012  {C1}
R501  3  N501  {R2}
L2  3  N015  {L1}
R54  3  N015  {Rs1}
L4  N015  N014  {L2}
R55  N015  N014  {Rs2}
L8  N013  N012  {L4}
R56  N013  N012  {Rs4}
L7  N009  N001  {L4}
R57  N009  N001  {Rs4}
L9  N001  N006  {L5}
R58  N001  N006  {Rs5}
C50  N001  N006  {C2}
L10  N012  N020  {L5}
R59  N012  N020  {Rs5}
C51  N012  N020  {C2}
R1  N002  1  {Rdc}
R6  N016  2  {Rdc}
R2  N006  N004  {dR6}
C1  N005  N004  {dC3}
L11  N008  N004  {dL3}
L12  N018  N019  {dL3}
C2  N008  N019  {ck}
R3  N006  N005  {dR5}
R4  N020  N022  {dR3}
C5  N022  N018  {dC3}
R5  N020  N018  {dR4}
L13  N006  N008  {dL3}
L14  N019  N020  {dL3}
R8  N004  N002  {dR6}
C6  N003  N002  {dC4}
L15  N007  N002  {dL4}
L16  N016  N017  {dL4}
C7  N007  N017  {ck}
R9  N004  N003  {dR5}
R10  N018  N021  {dR5}
C8  N021  N016  {dC4}
R11  N018  N016  {dR6}
L17  N004  N007  {dL4}
L18  N017  N018  {dL4}
K3  L5  L6  1
K2  L3  L4  1
K1  L1  L2  1
K4  L7  L8  1
K5  L9  L10  1
K6  L13  L14  L11  L12  0.9999
K7  L15  L16  L17  L18  0.9999
.ends  CMBNC
********
.subckt XS_7448010911_11m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.354999989271164
+  ck=9.15709522097963E-12
+  DC4=2.33921881864774E-10
+  DL4=1.09498807887576E-06
+  DR5=14846.5380859375
+  DR6=18534.806640625
+  DC3=3.33897409721118E-10
+  DL3=4.54652031578462E-08
+  DR3=1045.89575195313
+  DR4=88924.546875
+  L1=0.00869298074394464
+  L2=0.000467057310743257
+  L3=0.00135353673249483
+  L4=0.0000196324490389088
+  RS1=6607.99658203125
+  RS2=24180.732421875
+  RS3=9770.07421875
+  RS4=23873.265625
+  C1=4.78700456010839E-12
+  R2=3.01428484916687
+  C2=2.04170937934123E-08
+  L5=0.0000910909293452278
+  RS5=3.74318003654479
.ends XS_7448010911_11m
********
.subckt XS_7448011008_8m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.277999997138977
+  ck=6.0024012669968E-12
+  DC4=2.73229737446368E-11
+  DL4=8.14368092960649E-07
+  DR5=7221.44482421875
+  DR6=224451.9375
+  DC3=4.37110303508348E-09
+  DL3=5.67908315929344E-08
+  DR3=1169528.5
+  DR4=1024759.75
+  L1=0.0063436389900744
+  L2=0.00109203590545803
+  L3=0.000217066946788691
+  L4=0.00028052440029569
+  RS1=4582.064453125
+  RS2=7006.28369140625
+  RS3=47439.70703125
+  RS4=6601.64892578125
+  C1=3.50304941304502E-12
+  R2=2.29911279678345
+  C2=3.43900770491054E-13
+  L5=4.0811581891731E-10
+  RS5=0.41453218460083
.ends XS_7448011008_8m
********
.subckt XS_7448011305_5m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.168999999761581
+  ck=2.25999994678825E-14
+  DC4=3.65080535247309E-12
+  DL4=4.60730888107719E-07
+  DR5=3.52454352378845
+  DR6=6065.509765625
+  DC3=9.47457065060553E-13
+  DL3=2.40244109050991E-08
+  DR3=2051.99462890625
+  DR4=625860.9375
+  L1=0.00129573908634484
+  L2=0.00273191463202238
+  L3=0.000747762445826083
+  L4=0.000185409357072785
+  RS1=467.464172363281
+  RS2=2900.0927734375
+  RS3=5651.88671875
+  RS4=13813.4619140625
+  C1=3.34747615911291E-12
+  R2=1.03841233253479
+  C2=1.40755517050867E-13
+  L5=3.38628881879632E-11
+  RS5=2.2954523563385
.ends XS_7448011305_5m
********
.subckt XS_7448012002_1m6 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0860000029206276
+  ck=1.69815030093279E-12
+  DC4=1.18014398167027E-12
+  DL4=1.16388264359557E-07
+  DR5=61385.6328125
+  DR6=4105.31884765625
+  DC3=1.93209701709884E-11
+  DL3=6.56655041453291E-09
+  DR3=989.751708984375
+  DR4=2804660.25
+  L1=0.000852709752507508
+  L2=0.0000577403297938872
+  L3=0.000388926739105955
+  L4=0.000112803296360653
+  RS1=1605.56591796875
+  RS2=6322.48046875
+  RS3=88.5050964355469
+  RS4=1702.09875488281
+  C1=6.25561939488622E-13
+  R2=0.483416646718979
+  C2=6.73252102956212E-08
+  L5=0.0000249020140472567
+  RS5=42.8821487426758
.ends XS_7448012002_1m6
********
.subckt XS_7448012501_1m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.046000000089407
+  ck=1.64943427839737E-12
+  DC4=1.08074528544397E-16
+  DL4=9.4963432673012E-08
+  DR5=0.0133064752444625
+  DR6=3555.86938476563
+  DC3=5.14609996664903E-15
+  DL3=4.60131088786397E-09
+  DR3=0.0543990135192871
+  DR4=759.391662597656
+  L1=0.000334763084538281
+  L2=0.000046876710257493
+  L3=9.42685255722608E-06
+  L4=1.71062623621765E-07
+  RS1=366.980529785156
+  RS2=800.131530761719
+  RS3=1728.64892578125
+  RS4=12222.5107421875
+  C1=5.7560862543396E-13
+  R2=1.7486914396286
+  C2=1.55494833588982E-12
+  L5=0.00108504469972104
+  RS5=0.578695297241211
.ends XS_7448012501_1m
********
.subckt XS_7448013501_0m5 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0280000008642673
+  ck=1.49062598202299E-12
+  DC4=3.27661922388481E-14
+  DL4=5.61172690538569E-08
+  DR5=0.0279833115637302
+  DR6=2767.52563476563
+  DC3=1.85868383401414E-13
+  DL3=3.45350348318618E-09
+  DR3=9.8975133895874
+  DR4=660.719970703125
+  L1=0.000502295675687492
+  L2=0.000081971287727356
+  L3=1.63714980772056E-06
+  L4=0.0000160957752086688
+  RS1=516.5498046875
+  RS2=1053.02941894531
+  RS3=817.908447265625
+  RS4=2101.67431640625
+  C1=6.00873409188629E-13
+  R2=0.37173655629158
+  C2=4.61719800171068E-08
+  L5=0.0000011568936315598
+  RS5=0.534857392311096
.ends XS_7448013501_0m5
********
.subckt XS_7448014501_0m4 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0280000008642673
+  ck=4.0635138483236E-13
+  DC4=1.10570688889589E-12
+  DL4=3.89507022191538E-08
+  DR5=0.0495046675205231
+  DR6=2381.40185546875
+  DC3=2.40370576090956E-13
+  DL3=3.79364450964204E-09
+  DR3=1.26773536205292
+  DR4=14691058
+  L1=0.000311136245727539
+  L2=0.0000403032790927682
+  L3=2.99775706480432E-06
+  L4=8.61158605403034E-06
+  RS1=381.889678955078
+  RS2=724.102416992188
+  RS3=1262.0439453125
+  RS4=896.188537597656
+  C1=6.8501947820751E-13
+  R2=2.54812860488892
+  C2=3.12969011817543E-10
+  L5=0.000000796946153514
+  RS5=1.18781542778015
.ends XS_7448014501_0m4
********
.subckt M_7448030333_33m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0799999982118607
+  ck=1.73772524147964E-11
+  DC4=5.54359835813756E-10
+  DL4=1.26350835216726E-06
+  DR5=385153.40625
+  DR6=7327.30810546875
+  DC3=1.13417142344474E-09
+  DL3=4.8234202409958E-08
+  DR3=34255.38671875
+  DR4=22879832
+  L1=0.0247995257377625
+  L2=0.00917641445994377
+  L3=0.000879100640304387
+  L4=0.00202385382726789
+  RS1=4350.64990234375
+  RS2=7612.5126953125
+  RS3=2848405.25
+  RS4=9349.84765625
+  C1=8.26555230509785E-12
+  R2=37.8868217468262
+  C2=6.62411048324429E-06
+  L5=0.158110871911049
+  RS5=26937344
.ends M_7448030333_33m
********
.subckt M_7448030417_17m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0379999987781048
+  ck=1.562340014305E-11
+  DC4=3.28442655017636E-12
+  DL4=6.19997422290908E-07
+  DR5=46.389778137207
+  DR6=4362.0078125
+  DC3=1.29215174259241E-13
+  DL3=2.67301807355125E-08
+  DR3=100.374443054199
+  DR4=4953.90087890625
+  L1=0.0151557568460703
+  L2=0.00327215413562953
+  L3=0.000534946040716022
+  L4=0.000178101676283404
+  RS1=2870.03051757813
+  RS2=3019.1796875
+  RS3=6627.37109375
+  RS4=68425.8984375
+  C1=1.00611168701858E-11
+  R2=0.00632000016048551
+  C2=2.80000008638995E-13
+  L5=1.00000001335143E-10
+  RS5=1
.ends M_7448030417_17m
********
.subckt M_7448030509_9m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0219999998807907
+  ck=1.16532920466095E-11
+  DC4=5.88655253014325E-12
+  DL4=3.66745098290266E-07
+  DR5=125392.9609375
+  DR6=3499.224609375
+  DC3=1.43253794243625E-11
+  DL3=1.70972960233939E-08
+  DR3=5723.576171875
+  DR4=23600734208
+  L1=0.0120000001043081
+  L2=0.0020000000949949
+  L3=0.000500000023748726
+  L4=0.000150000007124618
+  RS1=1880
+  RS2=1900
+  RS3=4000
+  RS4=5000
+  C1=5.99999997602518E-12
+  R2=0.400000005960464
+  C2=2.80000008638995E-13
+  L5=1.00000001335143E-10
+  RS5=1
.ends M_7448030509_9m
********
.subckt M_7448031002_2m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00499999988824129
+  ck=2.87433163208284E-12
+  DC4=2.24046193923744E-12
+  DL4=5.47510552451058E-08
+  DR5=6099.224609375
+  DR6=3090.13427734375
+  DC3=1.15601473706095E-12
+  DL3=3.14217163399633E-09
+  DR3=845.783081054688
+  DR4=1123.61694335938
+  L1=0.00150000001303852
+  L2=0.000199999994947575
+  L3=0.0000599999984842725
+  L4=3.80000005861802E-06
+  RS1=400
+  RS2=500
+  RS3=1400
+  RS4=2300
+  C1=9.00000018087821E-13
+  R2=0.400000005960464
+  C2=2.80000008638995E-13
+  L5=1.00000001335143E-10
+  RS5=1
.ends M_7448031002_2m
********
.subckt M_7448031501_1m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0020000000949949
+  ck=2.57202570873305E-12
+  DC4=9.20577524800292E-13
+  DL4=3.5461745540033E-08
+  DR5=3732.66748046875
+  DR6=3327.22192382813
+  DC3=4.05753745489831E-13
+  DL3=2.54755616602154E-09
+  DR3=43.6796455383301
+  DR4=2774.19946289063
+  L1=0.00102942250669003
+  L2=0.0000951876281760633
+  L3=0.000016293502994813
+  L4=8.00845043613663E-07
+  RS1=322.377105712891
+  RS2=490.611419677734
+  RS3=1189.74926757813
+  RS4=3580.23168945313
+  C1=8.14731420349657E-13
+  R2=0.567472815513611
+  C2=3.6251337760633E-13
+  L5=1.25527727101726E-10
+  RS5=1.34631204605103
.ends M_7448031501_1m
********
.subckt L_7448040382_82m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.135000005364418
+  ck=5.98668475904063E-11
+  DC4=2.36828053912577E-13
+  DL4=3.88230228054454E-06
+  DR5=674.824829101563
+  DR6=9586.4306640625
+  DC3=1.14751775789901E-11
+  DL3=1.91542204319717E-09
+  DR3=21.6521663665771
+  DR4=512807040
+  L1=0.0829947218298912
+  L2=0.0101475343108177
+  L3=0.000536222942173481
+  L4=0.000365290936315432
+  RS1=20239.140625
+  RS2=28361.994140625
+  RS3=40298.8671875
+  RS4=5075.22265625
+  C1=2.74228764696183E-11
+  R2=0.286605805158615
+  C2=1.52322865432097E-08
+  L5=1.36148946694448E-06
+  RS5=1.43727397918701
.ends L_7448040382_82m
********
.subckt L_7448040435_35m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0640000030398369
+  ck=3.41574164786085E-11
+  DC4=1.86840939855187E-13
+  DL4=1.59136141064664E-06
+  DR5=834.48291015625
+  DR6=8056.29541015625
+  DC3=3.03443589699803E-11
+  DL3=5.20691649519289E-12
+  DR3=18.1167163848877
+  DR4=766605248
+  L1=0.0434059202671051
+  L2=0.00645833602175117
+  L3=0.00101479911245406
+  L4=0.00159177230671048
+  RS1=6704.43017578125
+  RS2=8743.3896484375
+  RS3=85064.4453125
+  RS4=9577.373046875
+  C1=1.56000004580825E-11
+  R2=0.104000002145767
+  C2=6.16184820501076E-07
+  L5=0.000372471375158057
+  RS5=302.954345703125
.ends L_7448040435_35m
********
.subckt L_7448040515_15m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0299999993294477
+  ck=2.09951552671006E-11
+  DC4=5.35570069196134E-13
+  DL4=6.62409661345009E-07
+  DR5=177.84440612793
+  DR6=5423.15185546875
+  DC3=2.21240335079864E-11
+  DL3=2.08324335559951E-09
+  DR3=25.7555999755859
+  DR4=790799680
+  L1=0.0313526727259159
+  L2=0.000232258913456462
+  L3=0.00022412148246076
+  L4=0.00299568800255656
+  RS1=2645.89135742188
+  RS2=3905.26733398438
+  RS3=60462.76953125
+  RS4=7249.16162109375
+  C1=7.88850842287081E-12
+  R2=2.64605188369751
+  C2=2.70506433253104E-07
+  L5=7.29241946828552E-06
+  RS5=18.6724090576172
.ends L_7448040515_15m
********
.subckt L_7448040707_7m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0149999996647239
+  ck=1.90952613964013E-12
+  DC4=1.85547193928826E-12
+  DL4=2.65392174014778E-07
+  DR5=7.91325426101685
+  DR6=5166.0283203125
+  DC3=1.44351640016249E-11
+  DL3=1.07662325235514E-11
+  DR3=20.0794124603271
+  DR4=573485056
+  L1=0.00819584168493748
+  L2=0.000104253798781428
+  L3=0.000717621645890176
+  L4=0.0000629422720521688
+  RS1=1761.64501953125
+  RS2=10478.921875
+  RS3=3873.51904296875
+  RS4=243.744842529297
+  C1=1.1602503896882E-12
+  R2=0.516414642333984
+  C2=1.75105725475078E-08
+  L5=1.16033824326678E-07
+  RS5=3.20607089996338
.ends L_7448040707_7m
********
.subckt L_7448041104_4m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00600000005215406
+  ck=4.35271480317412E-12
+  DC4=1.22982657044246E-11
+  DL4=1.54030630028501E-07
+  DR5=93915.5234375
+  DR6=3881.001953125
+  DC3=1.73222519661564E-10
+  DL3=4.94894569769144E-09
+  DR3=7971.07861328125
+  DR4=4366635
+  L1=0.00809952709823847
+  L2=0.000668641470838338
+  L3=0.0000666780688334256
+  L4=6.14096097706351E-06
+  RS1=967.972229003906
+  RS2=2600.03564453125
+  RS3=4233.78271484375
+  RS4=2245.02856445313
+  C1=1.06666368446251E-12
+  R2=0.651606798171997
+  C2=7.86708866939989E-08
+  L5=0.0000273303194262553
+  RS5=72.0766448974609
.ends L_7448041104_4m
********
.subckt L_7448041502_2m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00300000002607703
+  ck=6.9133678816391E-12
+  DC4=6.34493915740997E-11
+  DL4=7.75969937194532E-08
+  DR5=3128.60888671875
+  DR6=39471.07421875
+  DC3=1.05417675185914E-13
+  DL3=2.37918595935582E-09
+  DR3=274.328552246094
+  DR4=217580.609375
+  L1=0.00251754769124091
+  L2=0.000312576012220234
+  L3=0.0000346227570844349
+  L4=0.0000161843363457592
+  RS1=388.493408203125
+  RS2=987.174682617188
+  RS3=915.368774414063
+  RS4=2395.36376953125
+  C1=9.77613064286065E-13
+  R2=0.805560827255249
+  C2=2.31705442593072E-13
+  L5=2.30107197185525E-10
+  RS5=1.80797374248505
.ends L_7448041502_2m
********
.subckt L_7448041801_1m5 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0020000000949949
+  ck=3.53989407231303E-12
+  DC4=5.1319879742313E-14
+  DL4=7.49445590031428E-08
+  DR5=0.180175602436066
+  DR6=2204.73461914063
+  DC3=1.54048421154712E-12
+  DL3=4.0160017533708E-09
+  DR3=4.79514217376708
+  DR4=1317.73986816406
+  L1=0.00288988836109638
+  L2=0.000365983025403693
+  L3=0.000186753182788379
+  L4=0.0000447224119852763
+  RS1=335.088470458984
+  RS2=270.503509521484
+  RS3=602.089050292969
+  RS4=2233.65698242188
+  C1=1.2156046568651E-12
+  R2=0.46083676815033
+  C2=6.94929056521687E-08
+  L5=1.52263805830444E-06
+  RS5=1.9443267583847
.ends L_7448041801_1m5
********
.subckt L_7448042001_1m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0020000000949949
+  ck=3.54854752353251E-12
+  DC4=4.14999997799641E-14
+  DL4=4.42646452825102E-08
+  DR5=66.5085525512695
+  DR6=1859.89624023438
+  DC3=5.74410988609178E-14
+  DL3=2.73839506625961E-09
+  DR3=149.318984985352
+  DR4=2838661
+  L1=0.00169906951487064
+  L2=0.000165815101354383
+  L3=0.0000243897702603135
+  L4=0.0000125612896226812
+  RS1=320.175964355469
+  RS2=535.458984375
+  RS3=377.848846435547
+  RS4=1364.71984863281
+  C1=9.1106137391217E-13
+  R2=0.665103912353516
+  C2=5.02737158569744E-08
+  L5=1.29639533952286E-06
+  RS5=1.57858121395111
.ends L_7448042001_1m
********
.subckt XL_7448050219_190m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.270000010728836
+  ck=1.23371704020304E-13
+  DC4=3.71604483295762E-11
+  DL4=0.0000128481315186946
+  DR5=178.67951965332
+  DR6=344187.3125
+  DC3=2.00057175686608E-11
+  DL3=2.56449358276845E-11
+  DR3=56.1910705566406
+  DR4=10705463
+  L1=0.0765414461493492
+  L2=0.102970354259014
+  L3=0.0401266478002071
+  L4=0.00139641796704382
+  RS1=9568.2236328125
+  RS2=22181.89453125
+  RS3=44593.328125
+  RS4=43461.74609375
+  C1=3.402876938563E-11
+  R2=1.27523076534271
+  C2=4.27454374118952E-08
+  L5=1.66677966717543E-06
+  RS5=3.19618940353394
.ends XL_7448050219_190m
********
.subckt XL_7448050490_90m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0900000035762787
+  ck=1.74373070236516E-12
+  DC4=2.11479150163951E-11
+  DL4=5.81994072490488E-06
+  DR5=20.3653221130371
+  DR6=16725.390625
+  DC3=4.20192353134397E-12
+  DL3=1.90801571875454E-07
+  DR3=0.840387582778931
+  DR4=23183.978515625
+  L1=0.0633048415184021
+  L2=0.0527161695063114
+  L3=0.00819597952067852
+  L4=0.000813116610515863
+  RS1=7977.4462890625
+  RS2=21052.81640625
+  RS3=34378.23828125
+  RS4=21288.916015625
+  C1=1.64609645358915E-11
+  R2=0.626191973686218
+  C2=2.81210930097586E-08
+  L5=1.18083221423149E-06
+  RS5=0.190767958760262
.ends XL_7448050490_90m
********
.subckt XL_7448050530_30m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0390000008046627
+  ck=2.78509385692738E-11
+  DC4=2.03024242925211E-13
+  DL4=1.95580855688604E-06
+  DR5=1
+  DR6=8138.7958984375
+  DC3=9.44529177093756E-12
+  DL3=1.24510735055594E-10
+  DR3=6.0740008354187
+  DR4=968572096
+  L1=0.0328281410038471
+  L2=0.00365898618474603
+  L3=0.00248376303352416
+  L4=0.000128349827718921
+  RS1=6471.7998046875
+  RS2=5428.32861328125
+  RS3=22317.498046875
+  RS4=4520.37890625
+  C1=1.15296400898801E-11
+  R2=0.2381861358881
+  C2=1.21399867936134E-08
+  L5=3.81026836748788E-07
+  RS5=0.376253843307495
.ends XL_7448050530_30m
********
.subckt XL_7448051012_12m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0130000002682209
+  ck=1.29404375669856E-12
+  DC4=4.20166375650344E-12
+  DL4=5.41214205895812E-07
+  DR5=20.7590198516846
+  DR6=7527.47265625
+  DC3=3.50737125974498E-12
+  DL3=2.78807057441099E-08
+  DR3=1.97621190547943
+  DR4=164737248
+  L1=0.0120416963472962
+  L2=0.000347881024936214
+  L3=0.00163540430366993
+  L4=0.000174639615579508
+  RS1=2931.60400390625
+  RS2=9359.2822265625
+  RS3=3876.35083007813
+  RS4=4537.236328125
+  C1=1.85642104987005E-12
+  R2=0.539597749710083
+  C2=4.17126173601901E-08
+  L5=1.18381808533741E-06
+  RS5=1.67514705657959
.ends XL_7448051012_12m
********
.subckt XL_7448051804_4m5 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0130000002682209
+  ck=2.97196208615125E-12
+  DC4=4.81861989545807E-12
+  DL4=1.26532995636808E-07
+  DR5=127.255516052246
+  DR6=4357.1591796875
+  DC3=1.48002392134396E-13
+  DL3=6.84395544681138E-08
+  DR3=197.913146972656
+  DR4=2891.45288085938
+  L1=0.00452137878164649
+  L2=0.000352744333213195
+  L3=0.0000765442819101736
+  L4=0.0000105745393739198
+  RS1=1277.31860351563
+  RS2=2638.7890625
+  RS3=3978.26245117188
+  RS4=5125.6875
+  C1=2.37914874433309E-12
+  R2=0.514503955841064
+  C2=1.71329492815175E-08
+  L5=1.84958048521366E-06
+  RS5=1.35451459884644
.ends XL_7448051804_4m5
********
.subckt XL_7448052303_3m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0020000000949949
+  ck=7.26791630351054E-12
+  DC4=4.80728391122343E-12
+  DL4=1.6081330045381E-07
+  DR5=5729.1328125
+  DR6=5042.890625
+  DC3=1.36911168166498E-11
+  DL3=4.67032634787756E-09
+  DR3=587.157775878906
+  DR4=343236.9375
+  L1=0.00362045993097126
+  L2=0.000298893282888457
+  L3=0.0000368153596355114
+  L4=0.0000126412960526068
+  RS1=818.961853027344
+  RS2=2084.45874023438
+  RS3=1956.18017578125
+  RS4=3705.36303710938
+  C1=2.2923399289887E-12
+  R2=1.01931715011597
+  C2=1.24323151773353E-09
+  L5=0.0000270433974947082
+  RS5=168.055801391602
.ends XL_7448052303_3m
********
.subckt XL_7448052502_2m5 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00100000004749745
+  ck=8.29554849292313E-13
+  DC4=5.57796829558921E-11
+  DL4=1.43946996544742E-08
+  DR5=179.459518432617
+  DR6=4292.69921875
+  DC3=1.32724040091681E-12
+  DL3=1.11804851599118E-07
+  DR3=19.6222877502441
+  DR4=314498368
+  L1=0.00263017346151173
+  L2=0.000105558763607405
+  L3=0.00042800308438018
+  L4=8.12618600321002E-06
+  RS1=506.157012939453
+  RS2=2328.259765625
+  RS3=739.272888183594
+  RS4=10990.73046875
+  C1=1.75593979460931E-12
+  R2=1.93624866008759
+  C2=8.57131610132456E-08
+  L5=1.50932783071767E-06
+  RS5=1.53144800662994
.ends XL_7448052502_2m5
********
.subckt XL_7448053201_0m9 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0007999999797903
+  ck=1.2583327392221E-12
+  DC4=4.28396727814029E-12
+  DL4=4.20275760859568E-08
+  DR5=14.1212711334229
+  DR6=2775.19506835938
+  DC3=1.25812283768151E-12
+  DL3=3.20948245757791E-09
+  DR3=3.85115766525269
+  DR4=75660016
+  L1=0.000637456309050322
+  L2=0.000282176537439227
+  L3=0.0000572315802855883
+  L4=8.29354667075677E-06
+  RS1=125.572998046875
+  RS2=288.548736572266
+  RS3=825.164855957031
+  RS4=1331.63842773438
+  C1=2.28750894094854E-12
+  R2=5.2646689414978
+  C2=9.61421654094297E-12
+  L5=6.94416075930349E-06
+  RS5=5.94270849227905
.ends XL_7448053201_0m9
********
.subckt XXL_7448060535_35m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0839999988675117
+  ck=4.96077831591002E-12
+  DC4=1.98334820789015E-11
+  DL4=4.59804095953587E-06
+  DR5=56.921085357666
+  DR6=16531.955078125
+  DC3=8.23022986568001E-12
+  DL3=7.6840516172183E-09
+  DR3=10.2092542648315
+  DR4=250876416
+  L1=0.0213536079972982
+  L2=0.00678884657099843
+  L3=0.00133800145704299
+  L4=0.00335024832747877
+  RS1=20953.0625
+  RS2=84818.890625
+  RS3=2855.02490234375
+  RS4=4198.51025390625
+  C1=1.84510011436156E-11
+  R2=0.82143372297287
+  C2=6.83071235130228E-08
+  L5=2.43707540903415E-06
+  RS5=3.06103205680847
.ends XXL_7448060535_35m
********
.subckt XXL_7448060620_20m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0839999988675117
+  ck=6.01277014289359E-12
+  DC4=2.21204807943076E-11
+  DL4=3.06558172269433E-06
+  DR5=64.8782348632813
+  DR6=16196.1728515625
+  DC3=5.84814271661904E-12
+  DL3=2.1627684088088E-09
+  DR3=9.9702091217041
+  DR4=221807968
+  L1=0.0094672292470932
+  L2=0.00699292682111263
+  L3=0.00153509667143226
+  L4=0.00171207438688725
+  RS1=8777.9384765625
+  RS2=48527.07421875
+  RS3=868.967224121094
+  RS4=2137.66088867188
+  C1=1.78616791496333E-11
+  R2=0.608646094799042
+  C2=2.94578068604778E-08
+  L5=1.20935953873413E-06
+  RS5=1.22790324687958
.ends XXL_7448060620_20m
********
.subckt XXL_7448060814_14m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0189999993890524
+  ck=2.93837593146051E-11
+  DC4=2.35259562941792E-08
+  DL4=1.98842303689162E-06
+  DR5=5169.552734375
+  DR6=61153.6484375
+  DC3=2.04652362222578E-13
+  DL3=7.74112933754623E-08
+  DR3=640.601013183594
+  DR4=870.611022949219
+  L1=0.00970976520329714
+  L2=0.0021861451677978
+  L3=0.00137306982651353
+  L4=0.000958601187448949
+  RS1=9313.65234375
+  RS2=39263.6171875
+  RS3=1550.61120605469
+  RS4=3058.95092773438
+  C1=1.05860155710791E-11
+  R2=0.815732479095458
+  C2=4.0503952192239E-08
+  L5=0.000001271036126127
+  RS5=1.93002426624298
.ends XXL_7448060814_14m
********
.subckt XXL_7448061309_9m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00999999977648258
+  ck=4.06722919232827E-11
+  DC4=9.56819845576717E-10
+  DL4=1.31716421947203E-06
+  DR5=5652.556640625
+  DR6=7768.02001953125
+  DC3=3.17585888143235E-12
+  DL3=6.4419936052218E-08
+  DR3=412.457611083984
+  DR4=28079.703125
+  L1=0.00698916474357247
+  L2=0.00125871121417731
+  L3=0.00168122875038534
+  L4=0.00100450566969812
+  RS1=5720.06201171875
+  RS2=84753.640625
+  RS3=1992.466796875
+  RS4=4123.216796875
+  C1=1.80235514013471E-11
+  R2=1.04356241226196
+  C2=6.42019486463141E-08
+  L5=1.81636323759449E-06
+  RS5=2.22242593765259
.ends XXL_7448061309_9m
********
.subckt XXL_7448061507_7m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00600000005215406
+  ck=1.01505988944067E-12
+  DC4=1.75113951117467E-11
+  DL4=8.6810319999131E-07
+  DR5=10.5465259552002
+  DR6=4638.55908203125
+  DC3=2.46688300077061E-14
+  DL3=7.08466174614841E-08
+  DR3=0.705563604831696
+  DR4=10381737
+  L1=0.00506870495155454
+  L2=0.000874682678841054
+  L3=0.001658228575252
+  L4=0.000639679667074233
+  RS1=4715.02490234375
+  RS2=81134.6484375
+  RS3=1441.15991210938
+  RS4=3041.09594726563
+  C1=1.54103171196018E-11
+  R2=0.507139205932617
+  C2=3.47771305087008E-08
+  L5=8.98760902146023E-07
+  RS5=0.978153824806213
.ends XXL_7448061507_7m
********
.subckt XXL_7448062105_5m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00400000018998981
+  ck=2.95758348367592E-11
+  DC4=1.89999993277686E-14
+  DL4=6.64122239868448E-07
+  DR5=361.794647216797
+  DR6=3127.68603515625
+  DC3=7.73666634229508E-12
+  DL3=2.58115697704397E-08
+  DR3=710.999084472656
+  DR4=20627.453125
+  L1=0.00311436993069947
+  L2=0.000626115943305194
+  L3=0.000886573339812458
+  L4=0.000768705387599766
+  RS1=2827.06518554688
+  RS2=56696.171875
+  RS3=1517.8466796875
+  RS4=2845.55834960938
+  C1=1.39394138592985E-11
+  R2=0.461454510688782
+  C2=2.40371633708492E-08
+  L5=1.36279641083092E-06
+  RS5=0.996920466423035
.ends XXL_7448062105_5m
********
.subckt XXL_7448062603_3m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00300000002607703
+  ck=3.01888652964877E-11
+  DC4=5.33317801813121E-13
+  DL4=4.35371049434252E-07
+  DR5=1458.11145019531
+  DR6=3074.376953125
+  DC3=1.59807948124646E-11
+  DL3=1.70473359872858E-08
+  DR3=1219.49731445313
+  DR4=137247.921875
+  L1=0.00224578683264554
+  L2=0.000199999994947575
+  L3=0.00104663299862295
+  L4=0.000203529634745792
+  RS1=1250.37756347656
+  RS2=2809.2333984375
+  RS3=2588.65380859375
+  RS4=5889.67919921875
+  C1=1.18381771399556E-11
+  R2=1.23012852668762
+  C2=5.88680322266555E-08
+  L5=3.70975021724007E-06
+  RS5=1.8262939453125
.ends XXL_7448062603_3m
********
.subckt XXL_7448063801_1m5 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0020000000949949
+  ck=2.9528837708348E-11
+  DC4=1.81107342664411E-12
+  DL4=1.52490713389852E-07
+  DR5=136.359634399414
+  DR6=1262.17468261719
+  DC3=2.40683558153099E-12
+  DL3=8.66488214512628E-09
+  DR3=143.967742919922
+  DR4=609.906372070313
+  L1=0.000600735598709434
+  L2=0.00102119834627956
+  L3=0.000730740721337497
+  L4=0.000193675368791446
+  RS1=6
+  RS2=517.475830078125
+  RS3=1116.78527832031
+  RS4=4681.90576171875
+  C1=1.46737066941682E-11
+  R2=0.624236047267914
+  C2=3.67227634967549E-08
+  L5=1.21822552046069E-06
+  RS5=0.940431714057922
.ends XXL_7448063801_1m5
********
.subckt S_7448020680_80m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=1
+  ck=2.3668475904063E-11
+  DC4=1.706828053912577E-13
+  DL4=4.698230228054454E-06
+  DR5=674.824829101563
+  DR6=11886.4306640625
+  DC3=1.04751775789901E-12
+  DL3=1.91542204319717E-09
+  DR3=21.6521663665771
+  DR4=512807040
+  L1=0.08729947218298912
+  L2=0.0101475343108177
+  L3=0.000536222942173481
+  L4=0.000365290936315432
+  RS1=50239.140625
+  RS2=55361.994140625
+  RS3=40298.8671875
+  RS4=5075.22265625
+  C1=1.00810228764696183E-11
+  R2=28.6605805158615
+  C2=1.52322865432097E-08
+  L5=1.36148946694448E-06
+  RS5=1.43727397918701
.ends S_7448020680_80m
********
.subckt S_7448021230_30m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.28640000030398369
+  ck=2.01574164786085E-11
+  DC4=1.86840939855187E-13
+  DL4=1.59136141064664E-06
+  DR5=704.48291015625
+  DR6=6556.29541015625
+  DC3=3.03443589699803E-11
+  DL3=5.20691649519289E-12
+  DR3=18.1167163848877
+  DR4=766605248
+  L1=0.0208004059202671051
+  L2=0.00845833602175117
+  L3=0.00101479911245406
+  L4=0.00159177230671048
+  RS1=7904.43017578125
+  RS2=8743.3896484375
+  RS3=85064.4453125
+  RS4=19577.373046875
+  C1=0.92000004580825E-11
+  R2=0.104000002145767
+  C2=5.06184820501076E-07
+  L5=0.000372471375158057
+  RS5=302.954345703125
.ends S_7448021230_30m
********
.subckt S_7448022010_10m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.08509
+  ck=1.51552671006E-11
+  DC4=5.35570069196134E-13
+  DL4=6.62409661345009E-07
+  DR5=177.84440612793
+  DR6=3723.15185546875
+  DC3=2.21240335079864E-11
+  DL3=2.08324335559951E-09
+  DR3=25.7555999755859
+  DR4=790799680
+  L1=0.0082831352
+  L2=0.000232258913456462
+  L3=0.00022412148246076
+  L4=0.00299568800255656
+  RS1=2645.89135742188
+  RS2=3905.26733398438
+  RS3=60462.76953125
+  RS4=7249.16162109375
+  C1=7.88850842287081E-12
+  R2=2.64605188369751
+  C2=2.70506433253104E-07
+  L5=7.29241946828552E-06
+  RS5=18.6724090576172
.ends S_7448022010_10m
********
.subckt S_7448023005_5m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.040999996647239
+  ck=1.080952613964013E-12
+  DC4=1.85547193928826E-12
+  DL4=2.75392174014778E-07
+  DR5=7.91325426101685
+  DR6=3766.0283203125
+  DC3=1.44351640016249E-11
+  DL3=1.87662325235514E-11
+  DR3=20.0794124603271
+  DR4=573485056
+  L1=0.00519584168493748
+  L2=0.000204253798781428
+  L3=0.000717621645890176
+  L4=0.0000629422720521688
+  RS1=1561.64501953125
+  RS2=10478.921875
+  RS3=3173.51904296875
+  RS4=243.744842529297
+  C1=1.32802503896882E-12
+  R2=0.516414642333984
+  C2=1.75105725475078E-08
+  L5=1.16033824326678E-07
+  RS5=3.20607089996338
.ends S_7448023005_5m
********
.subckt S_7448024503_3m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0206
+  ck=3.900271480317412E-12
+  DC4=1.22982657044246E-11
+  DL4=1.54030630028501E-07
+  DR5=13915.5234375
+  DR6=3881.001953125
+  DC3=1.73222519661564E-10
+  DL3=4.94894569769144E-09
+  DR3=7971.07861328125
+  DR4=4366635
+  L1=0.002809952709823847
+  L2=0.0007168641470838338
+  L3=0.0000966780688334256
+  L4=6.14096097706351E-06
+  RS1=967.972229003906
+  RS2=2600.03564453125
+  RS3=4833.78271484375
+  RS4=2245.02856445313
+  C1=1.06666368446251E-12
+  R2=0.651606798171997
+  C2=5.86708866939989E-010
+  L5=0.0000273303194262553
+  RS5=72.0766448974609
.ends S_7448024503_3m
********
.subckt S_7448025003_2m5 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.00300000002607703
+  ck=4.5133678816391E-12
+  DC4=6.34493915740997E-11
+  DL4=13.15969937194532E-08
+  DR5=3128.60888671875
+  DR6=10471.07421875
+  DC3=2.05417675185914E-13
+  DL3=2.37918595935582E-09
+  DR3=274.328552246094
+  DR4=17580.609375
+  L1=0.0015502154769124091
+  L2=0.000812576012220234
+  L3=0.0001546227570844349
+  L4=0.0001061843363457592
+  RS1=388.493408203125
+  RS2=987.174682617188
+  RS3=915.368774414063
+  RS4=4195.36376953125
+  C1=9.97613064286065E-13
+  R2=0.805560827255249
+  C2=14.31705442593072E-14
+  L5=2.30107197185525E-10
+  RS5=1.80797374248505
.ends S_7448025003_2m5
********
.subckt S_7448026002_1m5 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0080000000949949
+  ck=3.23989407231303E-12
+  DC4=5.1319879742313E-16
+  DL4=7.69445590031428E-08
+  DR5=0.180175602436066
+  DR6=1754.73461914063
+  DC3=1.54048421154712E-16
+  DL3=4.0160017533708E-09
+  DR3=4.79514217376708
+  DR4=1317.73986816406
+  L1=0.00118988836109638
+  L2=0.0002305983025403693
+  L3=0.000206753182788379
+  L4=0.0000300147224119852763
+  RS1=335.088470458984
+  RS2=270.503509521484
+  RS3=602.089050292969
+  RS4=2833.65698242188
+  C1=1.0156046568651E-12
+  R2=0.46083676815033
+  C2=6.94929056521687E-08
+  L5=1.52263805830444E-06
+  RS5=1.9443267583847
.ends S_7448026002_1m5
********
.subckt S_7448027001_1m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0060000000949949
+  ck=3.4854752353251E-12
+  DC4=4.14999997799641E-14
+  DL4=5.1646452825102E-08
+  DR5=66.5085525512695
+  DR6=1249.89624023438
+  DC3=5.74410988609178E-14
+  DL3=2.73839506625961E-09
+  DR3=149.318984985352
+  DR4=2838661
+  L1=0.0009006951487064
+  L2=0.00025815101354383
+  L3=0.000050897702603135
+  L4=0.0000325612896226812
+  RS1=320.175964355469
+  RS2=535.458984375
+  RS3=377.848846435547
+  RS4=2064.71984863281
+  C1=1.1106137391217E-12
+  R2=0.665103912353516
+  C2=4.02737158569744E-08
+  L5=1.29639533952286E-06
+  RS5=1.57858121395111
.ends S_7448027001_1m
********
.subckt XL_7448051307_7m 1 2 3 4
X1  1  2  3  4  CMBNC  PARAMS:
+  Rdc=0.0130000002682209
+  ck=1.29404375669856E-12
+  DC4=6.80166375650344E-12
+  DL4=4.51214205895812E-07
+  DR5=1.7590198516846
+  DR6=3457.47265625
+  DC3=5.50737125974498E-12
+  DL3=2.78807057441099E-08
+  DR3=1.97621190547943
+  DR4=164737248
+  L1=0.0075416963472962
+  L2=0.000347881024936214
+  L3=0.00103540430366993
+  L4=0.000174639615579508
+  RS1=2931.60400390625
+  RS2=3059.2822265625
+  RS3=3576.35083007813
+  RS4=3537.236328125
+  C1=8.05642104987005E-12
+  R2=0.539597749710083
+  C2=4.17126173601901E-08
+  L5=1.18381808533741E-06
+  RS5=1.67514705657959
.ends XL_7448051307_7m
********