**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Polymer Capacitors
* Matchcode:             WCAP-PT5H
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 870235174001_390uF 1 2
Rser 1 3 0.00732480798856
Lser 2 4 3.866746561E-09
C1 3 4 0.00039
Rpar 3 4 12820.5128205128
.ends 870235174001_390uF
*******
.subckt 870235174002_470uF 1 2
Rser 1 3 0.00750285335959
Lser 2 4 4.014073535E-09
C1 3 4 0.00047
Rpar 3 4 10641.8918918919
.ends 870235174002_470uF
*******
.subckt 870235174003_560uF 1 2
Rser 1 3 0.00758797014666
Lser 2 4 6.337633943E-09
C1 3 4 0.00056
Rpar 3 4 8928.57142857143
.ends 870235174003_560uF
*******
.subckt 870235174004_680uF 1 2
Rser 1 3 0.00645535430737
Lser 2 4 5.020472116E-09
C1 3 4 0.00068
Rpar 3 4 14719.6261682243
.ends 870235174004_680uF
*******
.subckt 870235174005_820uF 1 2
Rser 1 3 0.00592887834629
Lser 2 4 5.12730135E-09
C1 3 4 0.00082
Rpar 3 4 12195.1219512195
.ends 870235174005_820uF
*******
.subckt 870235175006_1mF 1 2
Rser 1 3 0.00665519987306
Lser 2 4 4.759634087E-09
C1 3 4 0.001
Rpar 3 4 10000
.ends 870235175006_1mF
*******
.subckt 870235175007_1.2mF 1 2
Rser 1 3 0.00636308234344
Lser 2 4 4.906453052E-09
C1 3 4 0.0012
Rpar 3 4 8333.33333333333
.ends 870235175007_1.2mF
*******
.subckt 870235175008_1.5mF 1 2
Rser 1 3 0.0073612614271
Lser 2 4 7.253554609E-09
C1 3 4 0.0015
Rpar 3 4 6666.66666666667
.ends 870235175008_1.5mF
*******
.subckt 870235175009_2mF 1 2
Rser 1 3 0.00813172272965
Lser 2 4 4.08982236E-09
C1 3 4 0.002
Rpar 3 4 5000
.ends 870235175009_2mF
*******
.subckt 870235373001_100uF 1 2
Rser 1 3 0.00961672026554
Lser 2 4 3.675716308E-09
C1 3 4 0.0001
Rpar 3 4 100000
.ends 870235373001_100uF
*******
.subckt 870235373002_180uF 1 2
Rser 1 3 0.008655666397
Lser 2 4 5.241883503E-09
C1 3 4 0.00018
Rpar 3 4 55555.5555555556
.ends 870235373002_180uF
*******
.subckt 870235374003_180uF 1 2
Rser 1 3 0.00907602894231
Lser 2 4 5.51686224E-09
C1 3 4 0.00018
Rpar 3 4 55555.5555555556
.ends 870235374003_180uF
*******
.subckt 870235374004_220uF 1 2
Rser 1 3 0.00984408982682
Lser 2 4 4.861922421E-09
C1 3 4 0.00022
Rpar 3 4 45454.5454545455
.ends 870235374004_220uF
*******
.subckt 870235374005_270uF 1 2
Rser 1 3 0.0105329004472
Lser 2 4 5.358860986E-09
C1 3 4 0.00027
Rpar 3 4 37037.037037037
.ends 870235374005_270uF
*******
.subckt 870235374006_330uF 1 2
Rser 1 3 0.00879608874196
Lser 2 4 5.516689362E-09
C1 3 4 0.00033
Rpar 3 4 30303.0303030303
.ends 870235374006_330uF
*******
.subckt 870235375007_390uF 1 2
Rser 1 3 0.00870937254466
Lser 2 4 8.004209242E-09
C1 3 4 0.00039
Rpar 3 4 25641.0256410256
.ends 870235375007_390uF
*******
.subckt 870235375008_470uF 1 2
Rser 1 3 0.0104643985493
Lser 2 4 8.367752215E-09
C1 3 4 0.00047
Rpar 3 4 21276.5957446809
.ends 870235375008_470uF
*******
.subckt 870235375009_560uF 1 2
Rser 1 3 0.00822447237026
Lser 2 4 6.109749821E-09
C1 3 4 0.00056
Rpar 3 4 17857.1428571429
.ends 870235375009_560uF
*******
.subckt 870235673001_22uF 1 2
Rser 1 3 0.017
Lser 2 4 2.821763577E-09
C1 3 4 0.000022
Rpar 3 4 116666.666666667
.ends 870235673001_22uF
*******
.subckt 870235674003_39uF 1 2
Rser 1 3 0.0137038534727
Lser 2 4 3.28252174E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 870235674003_39uF
*******
.subckt 870235674004_68uF 1 2
Rser 1 3 0.004320076711
Lser 2 4 9.348374844E-09
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 870235674004_68uF
*******
.subckt 870235674005_82uF 1 2
Rser 1 3 0.00853441619684
Lser 2 4 3.520819747E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 870235674005_82uF
*******
.subckt 870235675002_33uF 1 2
Rser 1 3 0.0102799313364
Lser 2 4 4.320076711E-09
C1 3 4 0.000033
Rpar 3 4 151515.151515152
.ends 870235675002_33uF
*******
.subckt 870235675006_120uF 1 2
Rser 1 3 0.00851926760768
Lser 2 4 6.926634219E-09
C1 3 4 0.00012
Rpar 3 4 41666.6666666667
.ends 870235675006_120uF
*******
.subckt 870235675007_150uF 1 2
Rser 1 3 0.00858688403028
Lser 2 4 4.63632431E-09
C1 3 4 0.00015
Rpar 3 4 33333.3333333333
.ends 870235675007_150uF
*******
