**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT White Top view Ceramic LED
* Matchcode:              WL-SWTC
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-03-02
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 3535_158353027  1  2
D1 1 2 led
.MODEL led D
+ IS=213.37E-15
+ N=3.6731
+ RS=.10593
+ IKF=1.6190E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ TT=5.0000E-9
.ends
*****
.subckt 3535_158353030  1  2
D1 1 2 led
.MODEL led D
+ IS=213.37E-15
+ N=3.6731
+ RS=.10593
+ IKF=1.6190E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ TT=5.0000E-9
.ends
*****
.subckt 3535_158353040  1  2
D1 1 2 led
.MODEL led D
+ IS=213.37E-15
+ N=3.6731
+ RS=.10593
+ IKF=1.6190E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ TT=5.0000E-9
.ends
*****
.subckt 3535_158353050  1  2
D1 1 2 led
.MODEL led D
+ IS=213.37E-15
+ N=3.6731
+ RS=.10593
+ IKF=1.6190E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ TT=5.0000E-9
.ends
*****
.subckt 3535_158353060  1  2
D1 1 2 led
.MODEL led D
+ IS=213.37E-15
+ N=3.6731
+ RS=.10593
+ IKF=1.6190E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ TT=5.0000E-9
.ends
*****