**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Common Mode Power Line Choke 
* Matchcode:              WE-CMB NiZn
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-26
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt COM_IND  1  2  3  4  PARAMS:
L5  N011  N010  {L3}  
R50  N011  N010  {Rs3}  
C3  N500  N001  {C1}  
R500  4  N500  {R2}  
L1  4  N012  {L1}  
R51  4  N012  {Rs1}  
L3  N012  N011  {L2}  
R52  N012  N011  {Rs2}  
L6  N015  N014  {L3}  
R53  N015  N014  {Rs3}  
C4  N501  N013  {C1}  
R501  3  N501  {R2}  
L2  3  N016  {L1}  
R54  3  N016  {Rs1}  
L4  N016  N015  {L2}  
R55  N016  N015  {Rs2}  
L8  N014  N013  {L4}  
R56  N014  N013  {Rs4}  
L7  N010  N001  {L4}  
R57  N010  N001  {Rs4}  
L9  N001  N007  {L5}  
R58  N001  N007  {Rs5}  
C50  N001  N007  {C2}
L10  N013  N022  {L5}  
R59  N013  N022  {Rs5}  
C51  N013  N022  {C2}
L11  N007  N006  {L6}  
R60  N007  N006  {Rs6}  
C52  N007  N006  {C3}
L12  N022  N021  {L6}  
R61  N022  N021  {Rs6}  
C53  N022  N021  {C3}
R1  N002  1  {Rdc}    
R2  N004  N002  {dR4}    
C1  N003  N002  {dC3}    
L17  N008  N002  {dL3}    
L18  N017  N018  {dL3}    
C2  N008  N018  {ck}    
R3  N004  N003  {dR3}    
R4  N019  N023  {dR3}    
C9  N023  N017  {dC3}    
R5  N019  N017  {dR4}    
L19  N004  N008  {dL3}    
L20  N018  N019  {dL3}    
R6  N017  2  {Rdc}    
R8  N006  N004  {dR6}    
C10  N005  N004  {dC4}    
L13  N009  N004  {dL4}    
L14  N019  N020  {dL4}    
C11  N009  N020  {ck}    
R9  N006  N005  {dR5}    
R10  N021  N024  {dR5}    
C12  N024  N019  {dC4}    
R11  N021  N019  {dR6}    
L15  N006  N009  {dL4}    
L16  N020  N021  {dL4}    
K3  L5  L6  1    
K2  L3  L4  1    
K1  L1  L2  1    
K4  L7  L8  1    
K5  L9  L10  1    
K6  L11  L12  1    
K8  L17  L18  L19  L20  0.9999
K7  L13  L14  L15  L16  0.9999
.ends  COM_IND
*****
.subckt CMBNiZN 1 2 3 4 PARAMS:
+ L3=130u
+ Rs3=700
+ C1=1.8p
+ R2=1
+ L5=77u
+ C2=44.1p
+ Rs5=830
+ Rs1=0.1k
+ Rs2=10
+ Rs4=1
+ Rdc=1m
+ L1=0.8p
+ L2=1p
+ L4=1p
+ dR5=100
+ ck=7.5p
+ dL4=2n
+ dL3=0.05u
+ dC3=10.1p
+ dC4=1.1p
+ dR3=2.5k
+ dR6=1.53k
+ dR4=0.2k
L5 N009 N008 {L3}
C3 N002 N001 {C1}
L1 4 N010 {L1}
L3 N010 N009 {L2}
L6 N015 N014 {L3}
C4 N024 N013 {C1}
L2 3 N016 {L1}
L4 N016 N015 {L2}
L8 N014 N013 {L4}
L7 N008 N001 {L4}
L9 N001 N007 {L5}
L10 N013 N021 {L5}
R1 N003 1 {Rdc}
R2 N005 N003 {dR4}
C1 N004 N003 {dC3}
L17 N011 N003 {dL3}
L18 N017 N018 {dL3}
C2 N011 N018 {ck}
R3 N005 N004 {dR3}
R4 N019 N022 {dR3}
C9 N022 N017 {dC3}
R5 N019 N017 {dR4}
L19 N005 N011 {dL3}
L20 N018 N019 {dL3}
R6 N017 2 {Rdc}
R8 N007 N005 {dR6}
C10 N006 N005 {dC4}
L13 N012 N005 {dL4}
L14 N019 N020 {dL4}
C11 N012 N020 {ck}
R9 N007 N006 {dR5}
R10 N021 N023 {dR5}
C12 N023 N019 {dC4}
R11 N021 N019 {dR6}
L15 N007 N012 {dL4}
L16 N020 N021 {dL4}
R7 N001 N007 {Rs5}
C5 N001 N007 {C2}
R12 N013 N021 {Rs5}
C6 N013 N021 {C2}
R13 N008 N001 {Rs4}
R14 N009 N008 {Rs3}
R15 N010 N009 {Rs2}
R16 4 N010 {Rs1}
R17 N014 N013 {Rs4}
R18 N015 N014 {Rs3}
R19 N016 N015 {Rs2}
R20 3 N016 {Rs1}
R21 4 N002 {R2}
R22 3 N024 {R2}
K3 L5 L6 1
K2 L3 L4 1
K1 L1 L2 1
K4 L7 L8 1
K5 L9  L10 1
K7 L17 L18 L19 L20 0.9999
K6 L13 L14 L15 L16 0.9999
.ends
****
.subckt COM_IND23  1  2  3  4  PARAMS:    
R_R9  N12325  3  {R2}          
R_R8  N13265  N13287  {Rs4}          
Kn_K6  L_L11  L_L12            
+  L_L13  L_L14  0.9999          
R_R3  N12571  N12583  {Rs3}          
R_R10  N13777  4  {R2}          
C_C10  N13029  N12821  {ck}          
R_R20  N13215  N13229  {dR4}          
L_L11  N12821  N12295  {dL4}          
R_R17  N12267  N12273  {dR3}          
L_L8  N13265  N13287  {L4}          
R_R7  N13287  N13305  {Rs3}          
L_L9  N12295  N12307  {L5}          
Kn_K4  L_L7  L_L8  1          
R_R2  N12583  N12599  {Rs2}          
Kn_K5  L_L9  L_L10  1          
R_R16  N13229  N13249  {dR6}          
Kn_K7  L_L15  L_L16            
+  L_L17  L_L18  0.9999          
C_C5  N12273  N12289  {dC4}          
L_L6  N13287  N13305  {L3}          
L_L7  N12307  N12571  {L4}          
R_R6  N13305  N13319  {Rs2}          
R_R21  1  N12257  {Rdc}          
Kn_K3  L_L5  L_L6  1          
L_L16  N12257  N12799  {dL3}          
C_C8  N13215  N13741  {dC3}          
L_L18  N13023  N13215  {dL3}          
R_R1  N12599  3  {Rs1}          
R_R13  N12289  N12295  {dR5}          
L_L4  N13305  N13319  {L2}          
L_L5  N12571  N12583  {L3}          
R_R15  N13755  N13249  {dR5}          
R_R5  N13319  4  {Rs1}          
R_R18  N12257  N12273  {dR4}          
Kn_K2  L_L3  L_L4  1          
R_R19  N13741  N13229  {dR3}          
L_L15  N12799  N12273  {dL3}          
L_L17  N13229  N13023  {dL3}          
L_L3  N12583  N12599  {L2}          
R_R11  N12295  N12307  {Rs5}          
L_L2  N13319  4  {L1}          
C_C4  N13249  N13265  {C2}          
L_L10  N13249  N13265  {L5}          
Kn_K1  L_L1  L_L2  1          
R_R14  N12273  N12295  {dR6}          
C_C6  N13229  N13755  {dC4}          
L_L12  N12273  N12821  {dL4}          
L_L14  N13029  N13229  {dL4}          
L_L1  N12599  3  {L1}          
C_C1  N12307  N12325  {C1}          
R_R12  N13249  N13265  {Rs5}          
C_C2  N13265  N13777  {C1}          
R_R22  2  N13215  {Rdc}          
C_C9  N13023  N12799  {ck}          
R_R4  N12307  N12571  {Rs4}          
C_C3  N12295  N12307  {C2}          
L_L13  N13249  N13029  {dL4}          
C_C7  N12257  N12267  {dC3}                        
.ends  COM_IND23      
*****
.subckt XS_744841330_30u 1 2 3 4
X1  1  2  3  4  COM_IND  PARAMS:
+  L1=0.00002389
+  L2=0.00000429
+  L3=0.000001
+  L4=0.000001
+  L5=0.00000002526
+  L6=0.00000001951
+  C1=0.0000000000008638
+  C2=0.00000000000173
+  C3=0.0000000000002182
+  RS1=2340
+  RS2=2506
+  RS3=2254
+  RS4=88
+  RS5=0.09
+  RS6=783
+  R2=0.054
+  DL3=0.0000001489
+  DC3=3.13E-23
+  DL4=0.00000000085255
+  DC4=0.00000000000002967
+  DR3=425
+  DR4=5517
+  DR5=127
+  DR6=164
+  Rdc=14.665m
+  ck=4pF
.ends XS_744841330_30u
*****
.subckt XS_744841210_0.1m 1 2 3 4
X1  1  2  3  4  COM_IND  PARAMS:
+  L1=0.00006594
+  L2=0.0000059
+  L3=0.00000232
+  L4=0.00000103
+  L5=0.00000000628
+  L6=0.00000001156
+  C1=0.000000000000887951
+  C2=0.00000000000362
+  C3=0.00000000000006055
+  RS1=8033
+  RS2=5161
+  RS3=7079
+  RS4=7651
+  RS5=372
+  RS6=858
+  R2=11
+  DL3=0.00000038
+  DC3=3.58E-25
+  DL4=0.00000000032782
+  DC4=0.00000000001881
+  DR3=31
+  DR4=15181
+  DR5=1
+  DR6=4000
+  Rdc=51m
+  ck=4pF
.ends XS_744841210_0.1m
*****
.subckt XS_744841247_47u 1 2 3 4
X1  1  2  3  4  COM_IND  PARAMS:
+  L1=0.00003889
+  L2=0.00000429
+  L3=0.000001
+  L4=0.000009
+  L5=0.00000001526
+  L6=0.00000000726
+  C1=0.0000000000008638
+  C2=0.00000000000000473
+  C3=0.00000000000000923
+  RS1=4540
+  RS2=2506
+  RS3=2254
+  RS4=288
+  RS5=300
+  RS6=80
+  R2=0.054
+  DL3=0.00000027
+  DC3=0.0000000000007
+  DL4=0.000000001551
+  DC4=0.000000000000163
+  DR3=0.48
+  DR4=11680
+  DR5=0.78
+  DR6=7066
+  Rdc=23.9m
+  ck=4pF
.ends XS_744841247_47u
*****
.subckt S_7448421016_16u 1 2 3 4
X1  1  2  3  4  COM_IND  PARAMS:
+  L1=5u
+  L2=5u
+  L3=3u
+  L4=1.9u
+  L5=8.1n
+  L6=8n
+  C1=1.0p
+  C2=1.05p
+  C3=1f
+  RS1=900
+  RS2=250
+  RS3=500
+  RS4=880
+  RS5=900
+  RS6=1100
+  R2=1.41
+  DL3=0.000000055
+  DC3=0.0000000000018
+  DL4=0.00000000051
+  DC4=0.00000000000053
+  DR3=0.48
+  DR4=2680
+  DR5=0.78
+  DR6=866
+  Rdc=2.7m
+  ck=4pF
.ends S_7448421016_16u
*****
.subckt S_744842565_65u 1 2 3 4
X1  1  2  3  4  COM_IND  PARAMS:
+  L1=0.00002089
+  L2=0.00001829
+  L3=0.000003
+  L4=0.000003
+  L5=0.0000000126
+  L6=0.00000001951
+  C1=0.0000000000011638
+  C2=0.00000000000063
+  C3=0.0000000000002182
+  RS1=2740
+  RS2=2506
+  RS3=3254
+  RS4=508
+  RS5=500
+  RS6=100
+  R2=0.054
+  DL3=0.00000021
+  DC3=0.0000000000017
+  DL4=0.00000000389
+  DC4=0.00000000000033
+  DR3=0.48
+  DR4=8680
+  DR5=0.1
+  DR6=1066
+  Rdc=13m
+  ck=4pF
.ends S_744842565_65u
*****
.subckt S_744842742_42u 1 2 3 4
X1  1  2  3  4  COM_IND  PARAMS:
+  L1=.024m
+  L2=.01m
+  L3=0.7u
+  L4=0.5u
+  L5=12.4n
+  L6=33.4n
+  C1=1p
+  C2=.55p
+  C3=.65f
+  Rs1=2k
+  Rs2=3.8k
+  RS3=1100
+  RS4=90
+  RS5=900
+  RS6=200
+  R2=1.41
+  DL3=0.00000013
+  DC3=0.0000000000015
+  DL4=0.0000000011
+  DC4=0.00000000000000173
+  DR3=0.21
+  DR4=6680
+  DR5=385
+  DR6=1990.66
+  Rdc=8.1m
+  ck=4pF
.ends S_744842742_42u
*****
.subckt S_744842932_32u 1 2 3 4
X1  1  2  3  4  COM_IND  PARAMS:
+  L1=0.00001089
+  L2=0.00001029
+  L3=0.000003
+  L4=0.000009
+  L5=0.0000000126
+  L6=0.00000001951
+  C1=0.0000000000011638
+  C2=0.00000000000063
+  C3=0.0000000000002182
+  RS1=340
+  RS2=306
+  RS3=1254
+  RS4=2808
+  RS5=500
+  RS6=100
+  R2=0.054
+  DL3=0.0000001
+  DC3=0.0000000000021
+  DL4=0.0000000005
+  DC4=0.00000000000233
+  DR3=0.48
+  DR4=5680
+  DR5=0.58
+  DR6=766
+  Rdc=5.5m
+  ck=4pF
.ends S_744842932_32u
*****
.subckt XS_744841414_14u 1 2 3 4
X1  1  2  3  4  COM_IND23  PARAMS:
+  L1=1.54u
+  L2=1.23u
+  L3=0.70u
+  L4=9.9u
+  L5=8n
+  C1=800.06f
+  C2=900.02f
+  RS1=666.63
+  RS2=678.77
+  RS3=666.33
+  RS4=740
+  RS5=336.33
+  R2=12
+  DL3=0.000000067
+  DL4=0.00000000085
+  DC3=0.0000000000003
+  DC4=0.000000000000000002
+  DR3=6
+  DR4=3101
+  DR5=10
+  DR6=350
+  Rdc=6.043m
+  ck=4pF
.ends XS_744841414_14u
*****
*****
.subckt S_744842311_0.11m 1 2 3 4
X1  1  2  3  4  COM_IND23  PARAMS:
+  L1=.06m
+  L2=.06m
+  L3=3u
+  L4=9u
+  L5=33.4n
+  C1=1p
+  C2=.65p
+  Rs1=6k
+  Rs2=6k
+  RS3=800
+  RS4=90
+  RS5=1600
+  R2=1.41
+  DL3=0.00000038
+  DC3=0.0000000000016
+  DL4=0.00000000111
+  DC4=0.00000000000433
+  DR3=0.48
+  DR4=11680
+  DR5=0.58
+  DR6=1066
+  Rdc=31m
+  ck=4pF
.ends S_744842311_0.11m
*****
.subckt S_744842632_32u  1 2 3 4
X1  1  2  3  4  CMBNiZN  PARAMS:
+ L3=15u
+ Rs3=1200
+ C1=6.8p
+ R2=0.1
+ L5=13.5u
+ C2=0.97p
+ Rs5=4200
+ Rs1=0.0001k
+ Rs2=10
+ Rs4=1
+ Rdc=1m
+ L1=1p
+ L2=1p
+ L4=1p
+ dR5=0.00001
+ ck=0.75p
+ dL4=20n
+ dL3=0.055u
+ dC3=1p
+ dC4=0.001p
+ dR3=3.2k
+ dR6=8k
+ dR4=3k
.ends
*****
.subckt S_744842816_16u  1 2 3 4
X1  1  2  3  4  CMBNiZN  PARAMS:
+ L3=13u
+ Rs3=750
+ C1=8p
+ R2=0.1
+ L5=7u
+ C2=0.95p
+ Rs5=2660
+ Rs1=0.1k
+ Rs2=10
+ Rs4=1
+ Rdc=1m
+ L1=1p
+ L2=1p
+ L4=1p
+ dR5=1
+ ck=1.05p
+ dL4=7n
+ dL3=0.042u
+ dC3=0.9p
+ dC4=0.1p
+ dR3=13.2k
+ dR6=2.2k
+ dR4=1.6k
.ends
****