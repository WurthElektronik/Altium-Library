**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMD Flat Wire High Current Inductor
* Matchcode:             WE-HCIA
* Library Type:          LTspice
* Version:               rev22b
* Created/modified by:   Ella
* Date and Time:         06/08/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1050_7843250072_0.72u 1 2
Rp 1 2 463.339
Cp 1 2 3.29p
Rs 1 N3 0.00126
L1 N3 2 0.721u
.ends 1050_7843250072_0.72u
*******
.subckt 1050_784325012_1.2u 1 2
Rp 1 2 653.501
Cp 1 2 4.043p
Rs 1 N3 0.00186
L1 N3 2 1.076u
.ends 1050_784325012_1.2u
*******
.subckt 1050_784325018_1.8u 1 2
Rp 1 2 967.647
Cp 1 2 4.175p
Rs 1 N3 0.003
L1 N3 2 1.666u
.ends 1050_784325018_1.8u
*******
.subckt 1050_784325024_2.4u 1 2
Rp 1 2 1345
Cp 1 2 3.582p
Rs 1 N3 0.0049
L1 N3 2 2.34u
.ends 1050_784325024_2.4u
*******
.subckt 1050_784325033_3.3u 1 2
Rp 1 2 1628
Cp 1 2 4.811p
Rs 1 N3 0.0052
L1 N3 2 3.052u
.ends 1050_784325033_3.3u
*******
.subckt 1050_784325042_4.2u 1 2
Rp 1 2 2023
Cp 1 2 5.103p
Rs 1 N3 0.0071
L1 N3 2 3.887u
.ends 1050_784325042_4.2u
*******
.subckt 1050_784325055_5.2u 1 2
Rp 1 2 2383
Cp 1 2 5.366p
Rs 1 N3 0.0086
L1 N3 2 4.812u
.ends 1050_784325055_5.2u
*******
.subckt 1050_784325065_6.5u 1 2
Rp 1 2 2843
Cp 1 2 5.988p
Rs 1 N3 0.0105
L1 N3 2 6.051u
.ends 1050_784325065_6.5u
*******
.subckt 1050_784325078_7.8u 1 2
Rp 1 2 3201
Cp 1 2 6.36p
Rs 1 N3 0.0131
L1 N3 2 7.486u
.ends 1050_784325078_7.8u
*******
.subckt 1050_784325100_10u 1 2
Rp 1 2 4339
Cp 1 2 5.969p
Rs 1 N3 0.021
L1 N3 2 9.57u
.ends 1050_784325100_10u
*******
.subckt 1050_784325160_16.7u 1 2
Rp 1 2 6090
Cp 1 2 5.682p
Rs 1 N3 0.0345
L1 N3 2 16.881u
.ends 1050_784325160_16.7u
*******
.subckt 7050_7843140047_0.47u 1 2
Rp 1 2 335
Cp 1 2 0.75p
Rs 1 N3 0.00135
L1 N3 2 0.392u
.ends 7050_7843140047_0.47u
*******
.subckt 7050_784314011_1.1u 1 2
Rp 1 2 624
Cp 1 2 1.172p
Rs 1 N3 0.00315
L1 N3 2 0.998u
.ends 7050_784314011_1.1u
*******
.subckt 7050_784314033_3.3u 1 2
Rp 1 2 1464
Cp 1 2 1.854p
Rs 1 N3 0.009
L1 N3 2 2.899u
.ends 7050_784314033_3.3u
*******
.subckt 7050_784314049_4.9u 1 2
Rp 1 2 2179
Cp 1 2 1.495p
Rs 1 N3 0.0145
L1 N3 2 4.13u
.ends 7050_784314049_4.9u
*******
.subckt 7050_784314065_6.5u 1 2
Rp 1 2 3060
Cp 1 2 1.686p
Rs 1 N3 0.0215
L1 N3 2 5.988u
.ends 7050_784314065_6.5u
*******
.subckt 7050_784314100_10u 1 2
Rp 1 2 3970
Cp 1 2 1.69p
Rs 1 N3 0.033
L1 N3 2 8.728u
.ends 7050_784314100_10u
*******

