**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT Wire Wound Inductor
* Matchcode:             WE-ASI
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/8/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt L_74458303_3m 1 2
Rp 1 2 230068
Cp 1 2 20.444p
Rs 1 N3 3.5
L1 N3 2 2967u
.ends L_74458303_3m
*******
.subckt L_74458304_4.7m 1 2
Rp 1 2 253202
Cp 1 2 21.053p
Rs 1 N3 4.8
L1 N3 2 4578u
.ends L_74458304_4.7m
*******
.subckt L_74458306_6m 1 2
Rp 1 2 240832
Cp 1 2 19.431p
Rs 1 N3 6
L1 N3 2 5848u
.ends L_74458306_6m
*******
.subckt L_74458308_8m 1 2
Rp 1 2 298029
Cp 1 2 19.392p
Rs 1 N3 8
L1 N3 2 7616u
.ends L_74458308_8m
*******
.subckt M_744776333_3m 1 2
Rp 1 2 270119
Cp 1 2 11.101p
Rs 1 N3 7
L1 N3 2 2750u
.ends M_744776333_3m
*******
.subckt M_744776347_4.7m 1 2
Rp 1 2 320215
Cp 1 2 14.484p
Rs 1 N3 12
L1 N3 2 4040u
.ends M_744776347_4.7m
*******
.subckt M_744776360_6m 1 2
Rp 1 2 283414
Cp 1 2 14.6p
Rs 1 N3 16.7
L1 N3 2 5457u
.ends M_744776360_6m
*******
.subckt M_744776381_8m 1 2
Rp 1 2 400065
Cp 1 2 13.9p
Rs 1 N3 16
L1 N3 2 7471u
.ends M_744776381_8m
*******
.subckt Sensor_744775330_3m 1 2
Rp 1 2 307727
Cp 1 2 10.6p
Rs 1 N3 10
L1 N3 2 2878u
.ends Sensor_744775330_3m
*******
.subckt Sensor_744775347_4.7m 1 2
Rp 1 2 512966
Cp 1 2 11.1p
Rs 1 N3 13.8
L1 N3 2 4612u
.ends Sensor_744775347_4.7m
*******
.subckt Sensor_744775360_6m 1 2
Rp 1 2 467985
Cp 1 2 12.3p
Rs 1 N3 18
L1 N3 2 5715u
.ends Sensor_744775360_6m
*******
.subckt Sensor_744775380_8m 1 2
Rp 1 2 534565
Cp 1 2 6.622p
Rs 1 N3 25
L1 N3 2 7814u
.ends Sensor_744775380_8m
*******
.subckt Sensor_744775318_18m 1 2
Rp 1 2 1664000
Cp 1 2 9.78p
Rs 1 N3 72
L1 N3 2 16154u
.ends Sensor_744775318_18m
*******
