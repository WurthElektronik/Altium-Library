**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Ultraviolet Top LED Waterclear
* Matchcode:              WL-SUTW
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-08
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 2835_153283367A212  1  2
D1 1 2 led
.MODEL led D
+ IS=165.26E-21
+ N=3.3483
+ RS=2.0879
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_153283387A212  1  2
D1 1 2 led
.MODEL led D
+ IS=10.000E-21
+ N=2.7635
+ RS=.8188
+ IKF=6.8628
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=5.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_153283397A212  1  2
D1 1 2 led
.MODEL led D
+ IS=10.000E-21
+ N=2.7635
+ RS=.81889
+ IKF=6.9719
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=5.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_153283407A212  1  2
D1 1 2 led
.MODEL led D
+ IS=10.000E-21
+ N=2.7635
+ RS=.81889
+ IKF=6.9719
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=5.00E-6
+ TT=5.0000E-9
.ends
******