**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Toroidal Double Power Choke
* Matchcode:              WE-DCT
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt SH_744851016_0.16u  1  2  3  4  PARAMS:
+  Cww=5.47p
+  Rp1=448.31
+  Cp1=2.69p
+  Lp1=0.15u
+  Rp2=448.31
+  Cp2=2.69p
+  Lp2=0.15u
+  RDC1=0.0034
+  RDC2=0.0034
+  K=0.790569415042095
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851027_0.27u  1  2  3  4  PARAMS:
+  Cww=5.69p
+  Rp1=484.21
+  Cp1=2.9p
+  Lp1=0.23u
+  Rp2=484.21
+  Cp2=2.9p
+  Lp2=0.23u
+  RDC1=0.004
+  RDC2=0.004
+  K=0.805076485899413
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851039_0.39u  1  2  3  4  PARAMS:
+  Cww=9.85p
+  Rp1=560.46
+  Cp1=3.58p
+  Lp1=0.34u
+  Rp2=560.46
+  Cp2=3.58p
+  Lp2=0.34u
+  RDC1=0.0047
+  RDC2=0.0047
+  K=0.847318545736323
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851100_1u  1  2  3  4  PARAMS:
+  Cww=26.77p
+  Rp1=979.21
+  Cp1=4.21p
+  Lp1=0.93u
+  Rp2=979.21
+  Cp2=4.21p
+  Lp2=0.93u
+  RDC1=0.0074
+  RDC2=0.0074
+  K=0.888819441731559
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851102_100u  1  2  3  4  PARAMS:
+  Cww=83.4p
+  Rp1=12038.43
+  Cp1=6.01p
+  Lp1=98.69u
+  Rp2=12038.43
+  Cp2=6.01p
+  Lp2=98.69u
+  RDC1=0.265
+  RDC2=0.265
+  K=0.989696923305312
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851220_2.2u  1  2  3  4  PARAMS:
+  Cww=24.5p
+  Rp1=957.02
+  Cp1=4.22p
+  Lp1=1.86u
+  Rp2=957.02
+  Cp2=4.22p
+  Lp2=1.86u
+  RDC1=0.0074
+  RDC2=0.0074
+  K=0.939051746081217
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851221_22u  1  2  3  4  PARAMS:
+  Cww=53.07p
+  Rp1=3820.23
+  Cp1=6.74p
+  Lp1=19.85u
+  Rp2=3820.23
+  Cp2=6.74p
+  Lp2=19.85u
+  RDC1=0.034
+  RDC2=0.034
+  K=0.983962305264698
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851330_3.3u  1  2  3  4  PARAMS:
+  Cww=27.7p
+  Rp1=1315.27
+  Cp1=5.25p
+  Lp1=2.82u
+  Rp2=1315.27
+  Cp2=5.25p
+  Lp2=2.82u
+  RDC1=0.009
+  RDC2=0.009
+  K=0.955050371509907
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851471_47u  1  2  3  4  PARAMS:
+  Cww=63.16p
+  Rp1=6139.47
+  Cp1=5.56p
+  Lp1=42.39u
+  Rp2=6139.47
+  Cp2=5.56p
+  Lp2=42.39u
+  RDC1=0.13
+  RDC2=0.13
+  K=0.988228589285319
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_7448510091_91n  1  2  3  4  PARAMS:
+  Cww=3.4p
+  Rp1=431.01
+  Cp1=2.17p
+  Lp1=0.075u
+  Rp2=431.01
+  Cp2=2.17p
+  Lp2=0.075u
+  RDC1=0.0028
+  RDC2=0.0028
+  K=0.671229804574745
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt SH_744851470_4.7u  1  2  3  4  PARAMS:
+  Cww=31.6p
+  Rp1=1745
+  Cp1=6.15p
+  Lp1=4.25u
+  Rp2=1756
+  Cp2=6.22p
+  Lp2=4.28u
+  RDC1=0.0103
+  RDC2=0.0103
+  K=0.963702964743452
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
