*
*
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************

.subckt 760390012	1  2  3  6  5  4	
.param RxLkg=164.45ohm			
.param Leakage=0.197uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	174.902uH	Rser=135mohm	
Lpri2	2a	3	174.902uH	Rser=135mohm	
Lsec1	6	5	202.959uH	Rser=145mohm	
Lsec2	5	4	202.959uH	Rser=145mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=10.25pf			
.param Cprm2=10.1pf			
.param Rdmp1=146087.2ohm			
.param Rdmp2=146087.2ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 760390013	1  2  3  6  5  4	
.param RxLkg=109.34ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	174.9uH	Rser=125mohm	
Lpri2	2a	3	174.9uH	Rser=125mohm	
Lsec1	6	5	501.183uH	Rser=175mohm	
Lsec2	5	4	501.183uH	Rser=175mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=23.9pf			
.param Cprm2=23.9pf			
.param Rdmp1=95670.29ohm			
.param Rdmp2=95670.29ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 760390014	1  2  3  6  5  4	
.param RxLkg=244.26ohm			
.param Leakage=0.365uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	174.818uH	Rser=135mohm	
Lpri2	2a	3	174.818uH	Rser=135mohm	
Lsec1	6	5	299.26uH	Rser=155mohm	
Lsec2	5	4	299.26uH	Rser=155mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=15.95pf			
.param Cprm2=15.95pf			
.param Rdmp1=117109.46ohm			
.param Rdmp2=117109.46ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 760390015	1  2  3  6  5  4	
.param RxLkg=139.75ohm			
.param Leakage=0.36uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	174.82uH	Rser=150mohm	
Lpri2	2a	3	174.82uH	Rser=150mohm	
Lsec1	6	5	700uH	Rser=260mohm	
Lsec2	5	4	700uH	Rser=260mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=47.4pf			
.param Cprm2=47.05pf			
.param Rdmp1=67933.96ohm			
.param Rdmp2=67933.96ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends	

.subckt 750313710	1  2  3  6  5  4	
.param RxLkg=147.49ohm			
.param Leakage=0.216uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	191.392uH	Rser=140mohm	
Lpri2	2a	3	191.392uH	Rser=140mohm	
Lsec1	6	5	290.083uH	Rser=169mohm	
Lsec2	5	4	290.083uH	Rser=169mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=14pf			
.param Cprm2=14pf			
.param Rdmp1=130759.82ohm			
.param Rdmp2=130759.82ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends
		
.subckt 750316769	1  2  3  6  5  4	
.param RxLkg=51.64ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	124.9uH	Rser=200mohm	
Lpri2	2a	3	124.9uH	Rser=200mohm	
Lsec1	6	5	1491.736uH	Rser=575mohm	
Lsec2	5	4	1491.736uH	Rser=575mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=150pf			
.param Cprm2=150pf			
.param Rdmp1=32275.15ohm			
.param Rdmp2=32275.15ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316770	1  2  3  6  5  4	
.param RxLkg=63.25ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	124.9uH	Rser=160mohm	
Lpri2	2a	3	124.9uH	Rser=160mohm	
Lsec1	6	5	1057.851uH	Rser=393mohm	
Lsec2	5	4	1057.851uH	Rser=393mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=100pf			
.param Cprm2=100pf			
.param Rdmp1=39528.3ohm			
.param Rdmp2=39528.3ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750317331	1  2  3  6  5  4	
.param RxLkg=538.96ohm			
.param Leakage=2.5uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	1628.75uH	Rser=550mohm	
Lpri2	2a	3	1628.75uH	Rser=550mohm	
Lsec1	6	5	434.214uH	Rser=325mohm	
Lsec2	5	4	434.214uH	Rser=325mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=16.5pf			
.param Cprm2=16.5pf			
.param Rdmp1=351399.26ohm			
.param Rdmp2=351399.26ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750317828	1  2  3  6  5  4	
.param RxLkg=821.44ohm			
.param Leakage=4uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	1898uH	Rser=550mohm	
Lpri2	2a	3	1898uH	Rser=550mohm	
Lsec1	6	5	96.878uH	Rser=100mohm	
Lsec2	5	4	96.878uH	Rser=100mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=15.6pf			
.param Cprm2=15.6pf			
.param Rdmp1=390183.29ohm			
.param Rdmp2=390183.29ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750317829	1  2  3  6  5  4	
.param RxLkg=186.34ohm			
.param Leakage=0.6uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	719.7uH	Rser=400mohm	
Lpri2	2a	3	719.7uH	Rser=400mohm	
Lsec1	6	5	793.8uH	Rser=380mohm	
Lsec2	5	4	793.8uH	Rser=380mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=18pf			
.param Cprm2=18pf			
.param Rdmp1=223607ohm			
.param Rdmp2=223607ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750317830	1  2  3  6  5  4	
.param RxLkg=319.84ohm			
.param Leakage=0.8uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	849.6uH	Rser=350mohm	
Lpri2	2a	3	849.6uH	Rser=350mohm	
Lsec1	6	5	172.125uH	Rser=115mohm	
Lsec2	5	4	172.125uH	Rser=115mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=9.2pf			
.param Cprm2=9.2pf			
.param Rdmp1=339834.56ohm			
.param Rdmp2=339834.56ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750315225	1  2  3  6  5  4	
.param RxLkg=149.15ohm			
.param Leakage=0.145uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	96.928uH	Rser=73mohm	
Lpri2	2a	3	96.928uH	Rser=73mohm	
Lsec1	6	5	117.37uH	Rser=75mohm	
Lsec2	5	4	117.37uH	Rser=76mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=12.18pf			
.param Cprm2=12.18pf			
.param Rdmp1=99773.73ohm			
.param Rdmp2=99773.73ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750315226	1  2  3  6  5  4	
.param RxLkg=225.09ohm			
.param Leakage=0.253uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	96.874uH	Rser=73mohm	
Lpri2	2a	3	96.874uH	Rser=72mohm	
Lsec1	6	5	163.93uH	Rser=86mohm	
Lsec2	5	4	163.93uH	Rser=85mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=16.28pf			
.param Cprm2=16.28pf			
.param Rdmp1=86300.81ohm			
.param Rdmp2=86300.81ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750315227	1  2  3  6  5  4	
.param RxLkg=110.45ohm			
.param Leakage=0.155uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	96.923uH	Rser=75mohm	
Lpri2	2a	3	96.923uH	Rser=75mohm	
Lsec1	6	5	280.33uH	Rser=112mohm	
Lsec2	5	4	280.33uH	Rser=112mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=25.38pf			
.param Cprm2=25.38pf			
.param Rdmp1=69118.66ohm			
.param Rdmp2=69118.66ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750315228	1  2  3  6  5  4	
.param RxLkg=47009.44ohm			
.param Leakage=78.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	57.9uH	Rser=95mohm	
Lpri2	2a	3	57.9uH	Rser=94mohm	
Lsec1	6	5	388uH	Rser=204mohm	
Lsec2	5	4	388uH	Rser=203mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=35.66pf			
.param Cprm2=35.66pf			
.param Rdmp1=58310.94ohm			
.param Rdmp2=58310.94ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750314781	4  3  2  1  5  6  7  8	
.param RxLkg=848.95ohm			
.param Leakage=0.8uh			
Rlkg	4	4a	{RxLkg/2}	
L_Lkg	4	4a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	4a	3	39.6uH	Rser=43mohm	
Lpri2	2a	1	39.6uH	Rser=43mohm	
Lsec1	5	6	160uH	Rser=268mohm	
Lsec2	7	8	160uH	Rser=268mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=27.75pf			
.param Cprm2=27.75pf			
.param Rdmp1=42447.69ohm			
.param Rdmp2=42447.69ohm			
Cpri1	4	3	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	4	3	{Rdmp1}	
Rdmp2	2	1	{Rdmp2}	
Rg3	4	0	20meg	
Rg4	2	0	20meg	
Rg7	3	0	20meg	
Rg8	1	0	20meg	
Rg11	5	0	20meg	
Rg12	7	0	20meg	
Rg19	6	0	20meg	
Rg20	8	0	20meg	
.ends			

.subckt 750315213	3  2  1  6  7  8	
.param RxLkg=904.69ohm			
.param Leakage=1.95uh			
Rlkg	3	3a	{RxLkg/2}	
L_Lkg	3	3a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	3a	2	139.775uH	Rser=186mohm	
Lpri2	2a	1	139.775uH	Rser=188mohm	
Lsec1	6	7	140.75uH	Rser=275mohm	
Lsec2	7	8	140.75uH	Rser=279mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=41.26pf			
.param Cprm2=41.26pf			
.param Rdmp1=65300.13ohm			
.param Rdmp2=65300.13ohm			
Cpri1	3	2	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	3	2	{Rdmp1}	
Rdmp2	2	1	{Rdmp2}	
Rg3	3	0	20meg	
Rg7	2	0	20meg	
Rg8	1	0	20meg	
Rg11	6	0	20meg	
Rg19	7	0	20meg	
Rg20	8	0	20meg	
.ends			

.subckt 750315214	3  2  1  6  7  8	
.param RxLkg=1550.11ohm			
.param Leakage=2.61uh			
Rlkg	3	3a	{RxLkg/2}	
L_Lkg	3	3a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	3a	2	187.195uH	Rser=124mohm	
Lpri2	2a	1	187.195uH	Rser=126mohm	
Lsec1	6	7	11.781uH	Rser=38mohm	
Lsec2	7	8	11.781uH	Rser=39mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=18.8pf			
.param Cprm2=18.8pf			
.param Rdmp1=111952.38ohm			
.param Rdmp2=111952.38ohm			
Cpri1	3	2	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	3	2	{Rdmp1}	
Rdmp2	2	1	{Rdmp2}	
Rg3	3	0	20meg	
Rg7	2	0	20meg	
Rg8	1	0	20meg	
Rg11	6	0	20meg	
Rg19	7	0	20meg	
Rg20	8	0	20meg	
.ends	


.subckt 750315089	3  2  1  4  5  6	
.param RxLkg=434.51ohm			
.param Leakage=0.755uh			
Rlkg	3	3a	{RxLkg/2}	
L_Lkg	3	3a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	3a	2	169.623uH	Rser=874mohm	
Lpri2	2a	1	169.623uH	Rser=859mohm	
Lsec1	4	5	170uH	Rser=788mohm	
Lsec2	5	6	170uH	Rser=962mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=22.2pf			
.param Cprm2=22.2pf			
.param Rdmp1=97837.49ohm			
.param Rdmp2=97837.49ohm			
Cpri1	3	2	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	3	2	{Rdmp1}	
Rdmp2	2	1	{Rdmp2}	
Rg3	3	0	20meg	
Rg7	2	0	20meg	
Rg8	1	0	20meg	
Rg11	4	0	20meg	
Rg19	5	0	20meg	
Rg20	6	0	20meg	
.ends			

.subckt 750315090	3  2  1  4  5  6	
.param RxLkg=539.16ohm			
.param Leakage=0.4uh			
Rlkg	3	3a	{RxLkg/2}	
L_Lkg	3	3a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	3a	2	79.8uH	Rser=351mohm	
Lpri2	2a	1	79.8uH	Rser=348mohm	
Lsec1	4	5	80uH	Rser=243mohm	
Lsec2	5	6	80uH	Rser=303mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=8.6pf			
.param Cprm2=8.6pf			
.param Rdmp1=107832.53ohm			
.param Rdmp2=107832.53ohm			
Cpri1	3	2	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	3	2	{Rdmp1}	
Rdmp2	2	1	{Rdmp2}	
Rg3	3	0	20meg	
Rg7	2	0	20meg	
Rg8	1	0	20meg	
Rg11	4	0	20meg	
Rg19	5	0	20meg	
Rg20	6	0	20meg	
.ends			

.subckt 750315072	3  2  1  4  5  6	
.param RxLkg=498.17ohm			
.param Leakage=0.663uh			
Rlkg	3	3a	{RxLkg/2}	
L_Lkg	3	3a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	3a	2	204.669uH	Rser=687mohm	
Lpri2	2a	1	204.669uH	Rser=690mohm	
Lsec1	4	5	87.193uH	Rser=424mohm	
Lsec2	5	6	87.193uH	Rser=519mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=10.8pf			
.param Cprm2=10.8pf			
.param Rdmp1=154035.68ohm			
.param Rdmp2=154035.68ohm			
Cpri1	3	2	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	3	2	{Rdmp1}	
Rdmp2	2	1	{Rdmp2}	
Rg3	3	0	20meg	
Rg7	2	0	20meg	
Rg8	1	0	20meg	
Rg11	4	0	20meg	
Rg19	5	0	20meg	
Rg20	6	0	20meg	
.ends			


.subckt 750314706	3  2  1  4  5  6	
.param RxLkg=337.67ohm			
.param Leakage=0.438uh			
Rlkg	3	3a	{RxLkg/2}	
L_Lkg	3	3a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	3a	2	95.381uH	Rser=443mohm	
Lpri2	2a	1	95.381uH	Rser=447mohm	
Lsec1	4	5	309.744uH	Rser=714mohm	
Lsec2	5	6	309.744uH	Rser=880mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=22pf			
.param Cprm2=22pf			
.param Rdmp1=73700.72ohm			
.param Rdmp2=73700.72ohm			
Cpri1	3	2	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	3	2	{Rdmp1}	
Rdmp2	2	1	{Rdmp2}	
Rg3	3	0	20meg	
Rg7	2	0	20meg	
Rg8	1	0	20meg	
Rg11	4	0	20meg	
Rg19	5	0	20meg	
Rg20	6	0	20meg	
.ends			

.subckt 750311542	1  2  3  6  5  4	
.param RxLkg=408.25ohm			
.param Leakage=1uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	149.5uH	Rser=340mohm	
Lpri2	2a	3	149.5uH	Rser=340mohm	
Lsec1	6	5	1115.702uH	Rser=850mohm	
Lsec2	5	4	1115.702uH	Rser=850mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=50pf			
.param Cprm2=50pf			
.param Rdmp1=61237.49ohm			
.param Rdmp2=61237.49ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			


.subckt 750316853	1  2  3  6  5  4	
.param RxLkg=56.57ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	62.4uH	Rser=145mohm	
Lpri2	2a	3	62.4uH	Rser=145mohm	
Lsec1	6	5	1000uH	Rser=675mohm	
Lsec2	5	4	1000uH	Rser=675mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=250pf			
.param Cprm2=250pf			
.param Rdmp1=17677.74ohm			
.param Rdmp2=17677.74ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316854	1  2  3  6  5  4	
.param RxLkg=115.47ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	62.4uH	Rser=142.5mohm	
Lpri2	2a	3	62.4uH	Rser=142.5mohm	
Lsec1	6	5	390.625uH	Rser=425mohm	
Lsec2	5	4	390.625uH	Rser=425mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=60pf			
.param Cprm2=60pf			
.param Rdmp1=36084.33ohm			
.param Rdmp2=36084.33ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316855	1  2  3  6  5  4	
.param RxLkg=31.62ohm			
.param Leakage=0.25uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	62.375uH	Rser=225mohm	
Lpri2	2a	3	62.375uH	Rser=225mohm	
Lsec1	6	5	3062.5uH	Rser=2075mohm	
Lsec2	5	4	3062.5uH	Rser=2075mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=1250pf			
.param Cprm2=1250pf			
.param Rdmp1=7905.82ohm			
.param Rdmp2=7905.82ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316856	1  2  3  6  5  4	
.param RxLkg=44.72ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	62.4uH	Rser=147.5mohm	
Lpri2	2a	3	62.4uH	Rser=147.5mohm	
Lsec1	6	5	1361.111uH	Rser=1000mohm	
Lsec2	5	4	1361.111uH	Rser=1000mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=400pf			
.param Cprm2=400pf			
.param Rdmp1=13975.37ohm			
.param Rdmp2=13975.37ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316886	1  2  3  6  5  4	
.param RxLkg=319.21ohm			
.param Leakage=0.22uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	62.39uH	Rser=70mohm	
Lpri2	2a	3	62.39uH	Rser=70mohm	
Lsec1	6	5	85.069uH	Rser=88mohm	
Lsec2	5	4	85.069uH	Rser=88mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=9.5pf			
.param Cprm2=9.5pf			
.param Rdmp1=90684.43ohm			
.param Rdmp2=90684.43ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316887	1  2  3  6  5  4	
.param RxLkg=205.2ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	62.4uH	Rser=65mohm	
Lpri2	2a	3	62.4uH	Rser=65mohm	
Lsec1	6	5	173.611uH	Rser=188mohm	
Lsec2	5	4	173.611uH	Rser=188mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=19pf			
.param Cprm2=19pf			
.param Rdmp1=64123.83ohm			
.param Rdmp2=64123.83ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316888	1  2  3  6  5  4	
.param RxLkg=782.62ohm			
.param Leakage=0.35uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	62.325uH	Rser=90mohm	
Lpri2	2a	3	62.325uH	Rser=90mohm	
Lsec1	6	5	43.403uH	Rser=67.5mohm	
Lsec2	5	4	43.403uH	Rser=67.5mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=4pf			
.param Cprm2=4pf			
.param Rdmp1=139754.14ohm			
.param Rdmp2=139754.14ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750317072	1  2  3  6  5  4	
.param RxLkg=30.68ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	62.4uH	Rser=235mohm	
Lpri2	2a	3	62.4uH	Rser=235mohm	
Lsec1	6	5	2376.736uH	Rser=1725mohm	
Lsec2	5	4	2376.736uH	Rser=1725mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=850pf			
.param Cprm2=850pf			
.param Rdmp1=9586.96ohm			
.param Rdmp2=9586.96ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			



.subckt 750031160	3  2  1  4  5  6	
.param RxLkg=63.05ohm			
.param Leakage=0.28uh			
Rlkg	3	3a	{RxLkg/2}	
L_Lkg	3	3a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	3a	2	249.86uH	Rser=460mohm	
Lpri2	2a	1	249.86uH	Rser=460mohm	
Lsec1	4	5	1812.13uH	Rser=1200mohm	
Lsec2	5	6	1812.13uH	Rser=1200mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=98.6pf			
.param Cprm2=98.6pf			
.param Rdmp1=56297.34ohm			
.param Rdmp2=56297.34ohm			
Cpri1	3	2	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	3	2	{Rdmp1}	
Rdmp2	2	1	{Rdmp2}	
Rg3	3	0	20meg	
Rg7	2	0	20meg	
Rg8	1	0	20meg	
Rg11	4	0	20meg	
Rg19	5	0	20meg	
Rg20	6	0	20meg	
.ends			




.subckt 750316016	2  3  4  10  9  8  7  6	
.param RxLkg=696.31ohm			
.param Leakage=0.16uh			
Rlkg	2	2a	{RxLkg/2}	
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}	
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	3	21.92uH	Rser=54mohm	
Lpri2	3a	4	21.92uH	Rser=54mohm	
Lsec1	10	9	44.898uH	Rser=69mohm	
Lsec2	9	8	28.735uH	Rser=55mohm	
Lsec3	8	7	28.735uH	Rser=55mohm	
Lsec4	7	6	44.898uH	Rser=69mohm	
K Lpri1 Lpri2   Lsec1 Lsec2 Lsec3 Lsec4     1			
.param Cprm1=3pf			
.param Cprm2=3pf			
.param Rdmp1=95742.71ohm			
.param Rdmp2=95742.71ohm			
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	3	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}	
Rdmp2	3	4	{Rdmp2}	
Rg3	2	0	20meg	
Rg7	3	0	20meg	
Rg8	4	0	20meg	
Rg11	10	0	20meg	
Rg19	9	0	20meg	
Rg20	8	0	20meg	
Rg21	7	0	20meg	
Rg22	6	0	20meg	
.ends			

.subckt 750316017	2  3  4  10  9  8  7  6	
.param RxLkg=727.27ohm			
.param Leakage=0.16uh			
Rlkg	2	2a	{RxLkg/2}	
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}	
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	3	21.92uH	Rser=50mohm	
Lpri2	3a	4	21.92uH	Rser=50mohm	
Lsec1	10	9	64.653uH	Rser=120mohm	
Lsec2	9	8	16.163uH	Rser=44mohm	
Lsec3	8	7	16.163uH	Rser=44mohm	
Lsec4	7	6	64.653uH	Rser=120mohm	
K Lpri1 Lpri2   Lsec1 Lsec2 Lsec3 Lsec4     1			
.param Cprm1=2.75pf			
.param Cprm2=2.75pf			
.param Rdmp1=100000.06ohm			
.param Rdmp2=100000.06ohm			
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	3	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}	
Rdmp2	3	4	{Rdmp2}	
Rg3	2	0	20meg	
Rg7	3	0	20meg	
Rg8	4	0	20meg	
Rg11	10	0	20meg	
Rg19	9	0	20meg	
Rg20	8	0	20meg	
Rg21	7	0	20meg	
Rg22	6	0	20meg	
.ends			

.subckt 750316018	2  3  4  10  9  8  7  6	
.param RxLkg=603.02ohm			
.param Leakage=0.16uh			
Rlkg	2	2a	{RxLkg/2}	
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}	
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	3	21.92uH	Rser=51mohm	
Lpri2	3a	4	21.92uH	Rser=51mohm	
Lsec1	10	9	88uH	Rser=107mohm	
Lsec2	9	8	28.735uH	Rser=54mohm	
Lsec3	8	7	28.735uH	Rser=54mohm	
Lsec4	7	6	88uH	Rser=107mohm	
K Lpri1 Lpri2   Lsec1 Lsec2 Lsec3 Lsec4     1			
.param Cprm1=4pf			
.param Cprm2=4pf			
.param Rdmp1=82915.65ohm			
.param Rdmp2=82915.65ohm			
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	3	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}	
Rdmp2	3	4	{Rdmp2}	
Rg3	2	0	20meg	
Rg7	3	0	20meg	
Rg8	4	0	20meg	
Rg11	10	0	20meg	
Rg19	9	0	20meg	
Rg20	8	0	20meg	
Rg21	7	0	20meg	
Rg22	6	0	20meg	
.ends			

.subckt 750316019	2  3  4  10  9  8  7  6	
.param RxLkg=603.02ohm			
.param Leakage=0.16uh			
Rlkg	2	2a	{RxLkg/2}	
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}	
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	3	21.92uH	Rser=51mohm	
Lpri2	3a	4	21.92uH	Rser=51mohm	
Lsec1	10	9	88uH	Rser=107mohm	
Lsec2	9	8	28.735uH	Rser=54mohm	
Lsec3	8	7	28.735uH	Rser=54mohm	
Lsec4	7	6	88uH	Rser=107mohm	
K Lpri1 Lpri2   Lsec1 Lsec2 Lsec3 Lsec4     1			
.param Cprm1=4pf			
.param Cprm2=4pf			
.param Rdmp1=82915.65ohm			
.param Rdmp2=82915.65ohm			
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	3	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}	
Rdmp2	3	4	{Rdmp2}	
Rg3	2	0	20meg	
Rg7	3	0	20meg	
Rg8	4	0	20meg	
Rg11	10	0	20meg	
Rg19	9	0	20meg	
Rg20	8	0	20meg	
Rg21	7	0	20meg	
Rg22	6	0	20meg	
.ends			

.subckt 750316668	2  3  4  10  9  8  7  6	
.param RxLkg=696.31ohm			
.param Leakage=0.16uh			
Rlkg	2	2a	{RxLkg/2}	
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}	
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	3	21.92uH	Rser=54mohm	
Lpri2	3a	4	21.92uH	Rser=54mohm	
Lsec1	10	9	44.898uH	Rser=69mohm	
Lsec2	9	8	28.735uH	Rser=55mohm	
Lsec3	8	7	28.735uH	Rser=55mohm	
Lsec4	7	6	44.898uH	Rser=69mohm	
K Lpri1 Lpri2   Lsec1 Lsec2 Lsec3 Lsec4     1			
.param Cprm1=3pf			
.param Cprm2=3pf			
.param Rdmp1=95742.71ohm			
.param Rdmp2=95742.71ohm			
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	3	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}	
Rdmp2	3	4	{Rdmp2}	
Rg3	2	0	20meg	
Rg7	3	0	20meg	
Rg8	4	0	20meg	
Rg11	10	0	20meg	
Rg19	9	0	20meg	
Rg20	8	0	20meg	
Rg21	7	0	20meg	
Rg22	6	0	20meg	
.ends			

.subckt 750316669	2  3  4  10  9  8  7  6	
.param RxLkg=727.27ohm			
.param Leakage=0.16uh			
Rlkg	2	2a	{RxLkg/2}	
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}	
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	3	21.92uH	Rser=50mohm	
Lpri2	3a	4	21.92uH	Rser=50mohm	
Lsec1	10	9	64.653uH	Rser=120mohm	
Lsec2	9	8	16.163uH	Rser=44mohm	
Lsec3	8	7	16.163uH	Rser=44mohm	
Lsec4	7	6	64.653uH	Rser=120mohm	
K Lpri1 Lpri2   Lsec1 Lsec2 Lsec3 Lsec4     1			
.param Cprm1=2.75pf			
.param Cprm2=2.75pf			
.param Rdmp1=100000.06ohm			
.param Rdmp2=100000.06ohm			
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	3	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}	
Rdmp2	3	4	{Rdmp2}	
Rg3	2	0	20meg	
Rg7	3	0	20meg	
Rg8	4	0	20meg	
Rg11	10	0	20meg	
Rg19	9	0	20meg	
Rg20	8	0	20meg	
Rg21	7	0	20meg	
Rg22	6	0	20meg	
.ends			

.subckt 750316670	2  3  4  10  9  8  7  6	
.param RxLkg=603.02ohm			
.param Leakage=0.16uh			
Rlkg	2	2a	{RxLkg/2}	
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}	
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	3	21.92uH	Rser=51mohm	
Lpri2	3a	4	21.92uH	Rser=51mohm	
Lsec1	10	9	88uH	Rser=107mohm	
Lsec2	9	8	28.735uH	Rser=54mohm	
Lsec3	8	7	28.735uH	Rser=54mohm	
Lsec4	7	6	88uH	Rser=107mohm	
K Lpri1 Lpri2   Lsec1 Lsec2 Lsec3 Lsec4     1			
.param Cprm1=4pf			
.param Cprm2=4pf			
.param Rdmp1=82915.65ohm			
.param Rdmp2=82915.65ohm			
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	3	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}	
Rdmp2	3	4	{Rdmp2}	
Rg3	2	0	20meg	
Rg7	3	0	20meg	
Rg8	4	0	20meg	
Rg11	10	0	20meg	
Rg19	9	0	20meg	
Rg20	8	0	20meg	
Rg21	7	0	20meg	
Rg22	6	0	20meg	
.ends			

.subckt 750316671	2  3  4  10  9  8  7  6	
.param RxLkg=603.02ohm			
.param Leakage=0.16uh			
Rlkg	2	2a	{RxLkg/2}	
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}	
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	3	21.92uH	Rser=51mohm	
Lpri2	3a	4	21.92uH	Rser=51mohm	
Lsec1	10	9	88uH	Rser=107mohm	
Lsec2	9	8	28.735uH	Rser=54mohm	
Lsec3	8	7	28.735uH	Rser=54mohm	
Lsec4	7	6	88uH	Rser=107mohm	
K Lpri1 Lpri2   Lsec1 Lsec2 Lsec3 Lsec4     1			
.param Cprm1=4pf			
.param Cprm2=4pf			
.param Rdmp1=82915.65ohm			
.param Rdmp2=82915.65ohm			
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	3	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}	
Rdmp2	3	4	{Rdmp2}	
Rg3	2	0	20meg	
Rg7	3	0	20meg	
Rg8	4	0	20meg	
Rg11	10	0	20meg	
Rg19	9	0	20meg	
Rg20	8	0	20meg	
Rg21	7	0	20meg	
Rg22	6	0	20meg	
.ends	




.subckt 750315240	1  2  3  6  5  4	
.param RxLkg=532.24ohm			
.param Leakage=0.72uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	182.64uH	Rser=70mohm	
Lpri2	2a	3	182.64uH	Rser=70mohm	
Lsec1	6	5	225.926uH	Rser=62mohm	
Lsec2	5	4	225.926uH	Rser=62mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=12.5pf			
.param Cprm2=12.5pf			
.param Rdmp1=135277.82ohm			
.param Rdmp2=135277.82ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316031	1  2  3  6  5  4	
.param RxLkg=236.03ohm			
.param Leakage=0.38uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	119.81uH	Rser=64mohm	
Lpri2	2a	3	119.81uH	Rser=64mohm	
Lsec1	6	5	367.5uH	Rser=140mohm	
Lsec2	5	4	367.5uH	Rser=140mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=27pf			
.param Cprm2=27pf			
.param Rdmp1=74535.67ohm			
.param Rdmp2=74535.67ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316032	1  2  3  6  5  4	
.param RxLkg=198.95ohm			
.param Leakage=0.38uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	119.81uH	Rser=64mohm	
Lpri2	2a	3	119.81uH	Rser=64mohm	
Lsec1	6	5	480uH	Rser=160mohm	
Lsec2	5	4	480uH	Rser=160mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=38pf			
.param Cprm2=38pf			
.param Rdmp1=62827.83ohm			
.param Rdmp2=62827.83ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316033	1  2  3  6  5  4	
.param RxLkg=721.69ohm			
.param Leakage=0.5uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	119.75uH	Rser=64mohm	
Lpri2	2a	3	119.75uH	Rser=64mohm	
Lsec1	6	5	67.5uH	Rser=42mohm	
Lsec2	5	4	67.5uH	Rser=42mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=5pf			
.param Cprm2=5pf			
.param Rdmp1=173204.8ohm			
.param Rdmp2=173204.8ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			
		



.subckt 750313626	1  2  3  6  5  4	
.param RxLkg=139.17ohm			
.param Leakage=0.22uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	104.89uH	Rser=160mohm	
Lpri2	2a	3	104.89uH	Rser=160mohm	
Lsec1	6	5	420uH	Rser=225mohm	
Lsec2	5	4	420uH	Rser=225mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=29.75pf			
.param Cprm2=29.55pf			
.param Rdmp1=66421.41ohm			
.param Rdmp2=66421.41ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750313638	1  2  3  6  5  4	
.param RxLkg=340.21ohm			
.param Leakage=0.29uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	104.855uH	Rser=150mohm	
Lpri2	2a	3	104.855uH	Rser=150mohm	
Lsec1	6	5	186.667uH	Rser=150mohm	
Lsec2	5	4	186.667uH	Rser=150mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=8.65pf			
.param Cprm2=8.85pf			
.param Rdmp1=123180.34ohm			
.param Rdmp2=123180.34ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750313734	1  2  3  6  5  4	
.param RxLkg=475.5ohm			
.param Leakage=0.35uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	104.825uH	Rser=145mohm	
Lpri2	2a	3	104.825uH	Rser=145mohm	
Lsec1	6	5	129.63uH	Rser=130mohm	
Lsec2	5	4	129.63uH	Rser=130mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=6.45pf			
.param Cprm2=6.45pf			
.param Rdmp1=142649.1ohm			
.param Rdmp2=142649.1ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750313769	1  2  3  6  5  4	
.param RxLkg=214.31ohm			
.param Leakage=0.25uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	104.875uH	Rser=145mohm	
Lpri2	2a	3	104.875uH	Rser=145mohm	
Lsec1	6	5	291.667uH	Rser=185mohm	
Lsec2	5	4	291.667uH	Rser=185mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=16.2pf			
.param Cprm2=16.2pf			
.param Rdmp1=90010.21ohm			
.param Rdmp2=90010.21ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750343725	1  2  3  6  5  4	
.param RxLkg=97.29ohm			
.param Leakage=0.35uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	95.825uH	Rser=160mohm	
Lpri2	2a	3	95.825uH	Rser=160mohm	
Lsec1	6	5	1441.5uH	Rser=410mohm	
Lsec2	5	4	1441.5uH	Rser=410mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=168.5pf			
.param Cprm2=168.5pf			
.param Rdmp1=26686.15ohm			
.param Rdmp2=26686.15ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750342879	1  2  3  6  5  4	
.param RxLkg=121.97ohm			
.param Leakage=0.33uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	99.835uH	Rser=150mohm	
Lpri2	2a	3	99.835uH	Rser=150mohm	
Lsec1	6	5	1225uH	Rser=340mohm	
Lsec2	5	4	1225uH	Rser=340mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=91.5pf			
.param Cprm2=91.5pf			
.param Rdmp1=36960.84ohm			
.param Rdmp2=36960.84ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750343341	1  2  3  6  5  4	
.param RxLkg=149.4ohm			
.param Leakage=0.25uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	69.875uH	Rser=140mohm	
Lpri2	2a	3	69.875uH	Rser=140mohm	
Lsec1	6	5	462.857uH	Rser=230mohm	
Lsec2	5	4	462.857uH	Rser=230mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=50pf			
.param Cprm2=50pf			
.param Rdmp1=41832.88ohm			
.param Rdmp2=41832.88ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750315229	1  2  3  6  5  4	
.param RxLkg=226.87ohm			
.param Leakage=0.182uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	383.909uH	Rser=105mohm	
Lpri2	2a	3	383.909uH	Rser=105mohm	
Lsec1	6	5	303.407uH	Rser=114mohm	
Lsec2	5	4	303.407uH	Rser=114mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=2.095pf			
.param Cprm2=0pf			
.param Rdmp1=478661.7ohm			
.param Rdmp2=478661.7ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750315230	1  2  3  6  5  4	
.param RxLkg=168.19ohm			
.param Leakage=0.164uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	95.918uH	Rser=140mohm	
Lpri2	2a	3	95.918uH	Rser=141mohm	
Lsec1	6	5	50.777uH	Rser=161mohm	
Lsec2	5	4	50.777uH	Rser=161mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=12.38pf			
.param Cprm2=12.38pf			
.param Rdmp1=98453.19ohm			
.param Rdmp2=98453.19ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750315231	1  2  3  6  5  4	
.param RxLkg=237.3ohm			
.param Leakage=0.274uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	95.863uH	Rser=141mohm	
Lpri2	2a	3	95.863uH	Rser=140mohm	
Lsec1	6	5	36.355uH	Rser=161mohm	
Lsec2	5	4	36.355uH	Rser=161mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=17.36pf			
.param Cprm2=17.36pf			
.param Rdmp1=83141.32ohm			
.param Rdmp2=83141.32ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750315232	1  2  3  6  5  4	
.param RxLkg=125.99ohm			
.param Leakage=0.175uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	95.913uH	Rser=205mohm	
Lpri2	2a	3	95.913uH	Rser=205mohm	
Lsec1	6	5	24uH	Rser=175mohm	
Lsec2	5	4	24uH	Rser=175mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=25.12pf			
.param Cprm2=25.12pf			
.param Rdmp1=69116.65ohm			
.param Rdmp2=69116.65ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			



.subckt 750315371	1  2  3  6  5  4	
.param RxLkg=669.66ohm			
.param Leakage=0.255uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	24.873uH	Rser=25mohm	
Lpri2	2a	3	24.873uH	Rser=25mohm	
Lsec1	6	5	32.653uH	Rser=25mohm	
Lsec2	5	4	32.653uH	Rser=25mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=7.25pf			
.param Cprm2=7.25pf			
.param Rdmp1=65653.16ohm			
.param Rdmp2=65653.16ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316028	1  2  3  6  5  4	
.param RxLkg=205.06ohm			
.param Leakage=0.105uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	22.948uH	Rser=33mohm	
Lpri2	2a	3	22.948uH	Rser=33mohm	
Lsec1	6	5	67.592uH	Rser=48mohm	
Lsec2	5	4	67.592uH	Rser=48mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=14.25pf			
.param Cprm2=14.275pf			
.param Rdmp1=44917.03ohm			
.param Rdmp2=44917.03ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316029	1  2  3  6  5  4	
.param RxLkg=244.01ohm			
.param Leakage=0.157uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	22.922uH	Rser=33mohm	
Lpri2	2a	3	22.922uH	Rser=33mohm	
Lsec1	6	5	105.612uH	Rser=59mohm	
Lsec2	5	4	105.612uH	Rser=59mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=22.5pf			
.param Cprm2=23pf			
.param Rdmp1=35746.08ohm			
.param Rdmp2=35746.08ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316030	1  2  3  6  5  4	
.param RxLkg=539.82ohm			
.param Leakage=0.187uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	29.907uH	Rser=34mohm	
Lpri2	2a	3	29.907uH	Rser=34mohm	
Lsec1	6	5	16.875uH	Rser=28mohm	
Lsec2	5	4	16.875uH	Rser=28mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=5pf			
.param Cprm2=5pf			
.param Rdmp1=86602.59ohm			
.param Rdmp2=86602.59ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316818	1  2  3  6  5  4	
.param RxLkg=117.44ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	24.9uH	Rser=39mohm	
Lpri2	2a	3	24.9uH	Rser=39mohm	
Lsec1	6	5	306.25uH	Rser=220mohm	
Lsec2	5	4	306.25uH	Rser=220mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=145pf			
.param Cprm2=145pf			
.param Rdmp1=14680.51ohm			
.param Rdmp2=14680.51ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			

.subckt 750316819	1  2  3  6  5  4	
.param RxLkg=158.11ohm			
.param Leakage=0.2uh			
Rlkg	1	1a	{RxLkg/2}	
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}	
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	2	24.9uH	Rser=39mohm	
Lpri2	2a	3	24.9uH	Rser=39mohm	
Lsec1	6	5	206.641uH	Rser=175mohm	
Lsec2	5	4	206.641uH	Rser=175mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1			
.param Cprm1=80pf			
.param Cprm2=80pf			
.param Rdmp1=19764.23ohm			
.param Rdmp2=19764.23ohm			
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Cpri2	2	3	{Cprm2}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}	
Rdmp2	2	3	{Rdmp2}	
Rg3	1	0	20meg	
Rg7	2	0	20meg	
Rg8	3	0	20meg	
Rg11	6	0	20meg	
Rg19	5	0	20meg	
Rg20	4	0	20meg	
.ends			



