**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ATET
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 860130272001_47uF 1 2
Rser 1 3 0.95
Lser 2 4 0.000000003
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860130272001_47uF
*******
.subckt 860130273002_100uF 1 2
Rser 1 3 0.96297
Lser 2 4 7.731041053E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860130273002_100uF
*******
.subckt 860130274003_220uF 1 2
Rser 1 3 0.262
Lser 2 4 0.000000001
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860130274003_220uF
*******
.subckt 860130274004_330uF 1 2
Rser 1 3 0.23
Lser 2 4 0.0000000013
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860130274004_330uF
*******
.subckt 860130275005_470uF 1 2
Rser 1 3 0.205
Lser 2 4 0.000000002
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860130275005_470uF
*******
.subckt 860130275006_1mF 1 2
Rser 1 3 0.103
Lser 2 4 0.000000002
C1 3 4 0.001
Rpar 3 4 100000
.ends 860130275006_1mF
*******
.subckt 860130373001_33uF 1 2
Rser 1 3 1.19054473589
Lser 2 4 4.356034216E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860130373001_33uF
*******
.subckt 860130373002_47uF 1 2
Rser 1 3 0.65
Lser 2 4 5.100279947E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860130373002_47uF
*******
.subckt 860130373003_100uF 1 2
Rser 1 3 0.51
Lser 2 4 4.301638624E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860130373003_100uF
*******
.subckt 860130374004_220uF 1 2
Rser 1 3 0.222
Lser 2 4 0.000000002
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860130374004_220uF
*******
.subckt 860130375005_220uF 1 2
Rser 1 3 0.355
Lser 2 4 0.0000000011
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860130375005_220uF
*******
.subckt 860130375006_330uF 1 2
Rser 1 3 0.185
Lser 2 4 0.000000002
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860130375006_330uF
*******
.subckt 860130375007_470uF 1 2
Rser 1 3 0.153
Lser 2 4 0.000000002
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860130375007_470uF
*******
.subckt 860130375008_1mF 1 2
Rser 1 3 0.092
Lser 2 4 0.0000000035
C1 3 4 0.001
Rpar 3 4 100000
.ends 860130375008_1mF
*******
.subckt 860130378009_1mF 1 2
Rser 1 3 0.1
Lser 2 4 0.000000003
C1 3 4 0.001
Rpar 3 4 100000
.ends 860130378009_1mF
*******
.subckt 860130473001_22uF 1 2
Rser 1 3 0.55
Lser 2 4 4.075745866E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860130473001_22uF
*******
.subckt 860130473002_33uF 1 2
Rser 1 3 0.720217743803
Lser 2 4 5.300851003E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860130473002_33uF
*******
.subckt 860130473003_47uF 1 2
Rser 1 3 0.64
Lser 2 4 3.711513552E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860130473003_47uF
*******
.subckt 860130474004_100uF 1 2
Rser 1 3 0.275
Lser 2 4 0.0000000022
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860130474004_100uF
*******
.subckt 860130475005_100uF 1 2
Rser 1 3 0.27
Lser 2 4 7.038660156E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860130475005_100uF
*******
.subckt 860130475006_220uF 1 2
Rser 1 3 0.193
Lser 2 4 0.0000000017
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860130475006_220uF
*******
.subckt 860130475007_330uF 1 2
Rser 1 3 0.095
Lser 2 4 0.000000003
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860130475007_330uF
*******
.subckt 860130475008_470uF 1 2
Rser 1 3 0.081
Lser 2 4 0.000000004
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860130475008_470uF
*******
.subckt 860130478009_470uF 1 2
Rser 1 3 0.094
Lser 2 4 0.000000006
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860130478009_470uF
*******
.subckt 860130478010_1mF 1 2
Rser 1 3 0.062
Lser 2 4 0.000000014
C1 3 4 0.001
Rpar 3 4 100000
.ends 860130478010_1mF
*******
.subckt 860130573001_22uF 1 2
Rser 1 3 0.55
Lser 2 4 3.948129143E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 860130573001_22uF
*******
.subckt 860130574002_33uF 1 2
Rser 1 3 0.29
Lser 2 4 0.000000005
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860130574002_33uF
*******
.subckt 860130574003_47uF 1 2
Rser 1 3 0.34
Lser 2 4 4.550322687E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860130574003_47uF
*******
.subckt 860130575004_100uF 1 2
Rser 1 3 0.43
Lser 2 4 0.0000000008
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860130575004_100uF
*******
.subckt 860130575005_220uF 1 2
Rser 1 3 0.135
Lser 2 4 0.000000003
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860130575005_220uF
*******
.subckt 860130575006_330uF 1 2
Rser 1 3 0.097
Lser 2 4 0.000000005
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860130575006_330uF
*******
.subckt 860130578007_330uF 1 2
Rser 1 3 0.099
Lser 2 4 0.000000007
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860130578007_330uF
*******
.subckt 860130578008_470uF 1 2
Rser 1 3 0.074
Lser 2 4 0.000000007
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860130578008_470uF
*******
.subckt 860130580009_1mF 1 2
Rser 1 3 0.044
Lser 2 4 0.000000008
C1 3 4 0.001
Rpar 3 4 100000
.ends 860130580009_1mF
*******
.subckt 860130673001_10uF 1 2
Rser 1 3 0.6
Lser 2 4 3.698884681E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860130673001_10uF
*******
.subckt 860130673002_22uF 1 2
Rser 1 3 0.7
Lser 2 4 3.642276759E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860130673002_22uF
*******
.subckt 860130674003_33uF 1 2
Rser 1 3 0.29
Lser 2 4 0.0000000045
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860130674003_33uF
*******
.subckt 860130674004_47uF 1 2
Rser 1 3 0.45
Lser 2 4 4.6607845E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860130674004_47uF
*******
.subckt 860130675005_47uF 1 2
Rser 1 3 0.28
Lser 2 4 6.384870597E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860130675005_47uF
*******
.subckt 860130675006_100uF 1 2
Rser 1 3 0.212
Lser 2 4 0.0000000025
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860130675006_100uF
*******
.subckt 860130675007_220uF 1 2
Rser 1 3 0.131
Lser 2 4 0.0000000045
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860130675007_220uF
*******
.subckt 860130678008_220uF 1 2
Rser 1 3 0.105
Lser 2 4 0.0000000065
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860130678008_220uF
*******
.subckt 860130678009_330uF 1 2
Rser 1 3 0.082
Lser 2 4 0.000000007
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860130678009_330uF
*******
.subckt 860130678010_470uF 1 2
Rser 1 3 0.061
Lser 2 4 0.00000001
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860130678010_470uF
*******
.subckt 860130873001_470nF 1 2
Rser 1 3 0.9
Lser 2 4 3.689993692E-09
C1 3 4 0.00000047
Rpar 3 4 33333333.3333333
.ends 860130873001_470nF
*******
.subckt 860130873002_1uF 1 2
Rser 1 3 0.8
Lser 2 4 4.023385572E-09
C1 3 4 0.000001
Rpar 3 4 33333333.3333333
.ends 860130873002_1uF
*******
.subckt 860130873003_2.2uF 1 2
Rser 1 3 1.01490022899
Lser 2 4 3.580350161E-09
C1 3 4 0.0000022
Rpar 3 4 33333333.3333333
.ends 860130873003_2.2uF
*******
.subckt 860130873004_3.3uF 1 2
Rser 1 3 0.716082878235
Lser 2 4 3.861516865E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 860130873004_3.3uF
*******
.subckt 860130873005_4.7uF 1 2
Rser 1 3 1.0128660645
Lser 2 4 3.517981985E-09
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 860130873005_4.7uF
*******
.subckt 860130874006_10uF 1 2
Rser 1 3 0.37
Lser 2 4 5.573643346E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860130874006_10uF
*******
.subckt 860130875007_22uF 1 2
Rser 1 3 0.198436668232
Lser 2 4 6.325531422E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860130875007_22uF
*******
.subckt 860130875008_33uF 1 2
Rser 1 3 0.13
Lser 2 4 0.000000008
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860130875008_33uF
*******
.subckt 860130875009_47uF 1 2
Rser 1 3 0.105
Lser 2 4 0.00000001
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860130875009_47uF
*******
.subckt 860130878010_47uF 1 2
Rser 1 3 0.099
Lser 2 4 0.00000001
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860130878010_47uF
*******
.subckt 860130878011_100uF 1 2
Rser 1 3 0.063
Lser 2 4 0.0000000124
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860130878011_100uF
*******
.subckt 860131173001_1uF 1 2
Rser 1 3 1.86471696741
Lser 2 4 3.090425884E-09
C1 3 4 0.000001
Rpar 3 4 83333333.3333333
.ends 860131173001_1uF
*******
.subckt 860131173002_2.2uF 1 2
Rser 1 3 1.84349270446
Lser 2 4 3.530267079E-09
C1 3 4 0.0000022
Rpar 3 4 45454545.4545455
.ends 860131173002_2.2uF
*******
.subckt 860131174003_3.3uF 1 2
Rser 1 3 1.22264289826
Lser 2 4 3.436322371E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 860131174003_3.3uF
*******
.subckt 860131175004_4.7uF 1 2
Rser 1 3 1.12572119109
Lser 2 4 4.218792702E-09
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 860131175004_4.7uF
*******
.subckt 860131175005_10uF 1 2
Rser 1 3 0.815834470101
Lser 2 4 5.102550051E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860131175005_10uF
*******
.subckt 860131178006_22uF 1 2
Rser 1 3 0.538705989803
Lser 2 4 6.024415617E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860131178006_22uF
*******
.subckt 860131178007_33uF 1 2
Rser 1 3 0.366548331185
Lser 2 4 6.299102934E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860131178007_33uF
*******
.subckt 860131180008_47uF 1 2
Rser 1 3 0.18
Lser 2 4 8.98270434E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860131180008_47uF
*******
.subckt 860131274001_1uF 1 2
Rser 1 3 1.5065112609
Lser 2 4 3.837025608E-09
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 860131274001_1uF
*******
.subckt 860131274002_2.2uF 1 2
Rser 1 3 1.81673881249
Lser 2 4 7.183855007E-09
C1 3 4 0.0000022
Rpar 3 4 45454545.4545455
.ends 860131274002_2.2uF
*******
.subckt 860131275003_3.3uF 1 2
Rser 1 3 1.17092220856
Lser 2 4 4.136467848E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 860131275003_3.3uF
*******
.subckt 860131275004_4.7uF 1 2
Rser 1 3 1.01316567389
Lser 2 4 5.439895523E-09
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 860131275004_4.7uF
*******
.subckt 860131275005_10uF 1 2
Rser 1 3 0.721442464128
Lser 2 4 4.827049762E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860131275005_10uF
*******
.subckt 860131278006_10uF 1 2
Rser 1 3 0.580505434841
Lser 2 4 6.31541815E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860131278006_10uF
*******
.subckt 860131278007_22uF 1 2
Rser 1 3 0.578512003787
Lser 2 4 6.6242581E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860131278007_22uF
*******
.subckt 860131280008_33uF 1 2
Rser 1 3 0.493728689076
Lser 2 4 1.190214525E-08
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860131280008_33uF
*******
.subckt 860131280009_47uF 1 2
Rser 1 3 0.31
Lser 2 4 0.0000000003
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860131280009_47uF
*******
