**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Common Mode Power Line Choke (Horizontal)
* Matchcode:              WE-CMBH 
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Ella      
* Date and Time:          2022-07-19
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.SUBCKT L_744834101_1m  1  2  3  4
X1  1  2  3  4  CMBH  PARAMS:
+  L1=485.0122u
+  L2=321.4326u
+  L3=76.9226u
+  L4=1.2315u
+  L5=193.3875u
+  C1=19.0082p
+  C2=2.9783p
+  Rs1=2.5613k
+  Rs2=1.6990k
+  Rs3=3.7563k
+  Rs4=30.1669k
+  Rs5=3.0982k
+  R2=44.8612
+  dL3=318.6802n
+  dC3=5.7509p
+  dL4=11.9625n
+  dC4=5.4629p
+  dR3=479.4630m
+  dR4=438.6748
+  dR5=779.6469m
+  dR6=166.2752
+  Rdc=12.5m
+  ck=201.6390f
.ends  
**** 
.SUBCKT L_744834622_2.2m  1  2  3  4
X1  1  2  3  4  CMBH  PARAMS:
+  L1=2.4759m
+  L2=256.6851u
+  L3=13.1500u
+  L4=100.0003n
+  L5=169.9280n
+  C1=12.0967p
+  C2=100.0001f
+  Rs1=17.0959k
+  Rs2=2.0011k
+  Rs3=200.0031
+  Rs4=260.0000
+  Rs5=459.9999
+  R2=1.4100
+  dL3=848.8863n
+  dC3=5.0791p
+  dL4=13.6276n
+  dC4=13.8449p
+  dR3=490.0099m
+  dR4=5.8802k
+  dR5=16.9990
+  dR6=866.0010
+  Rdc=22m
+  ck=100f
.ends 
****
.SUBCKT L_744834433_3.3m  1  2  3  4
X1  1  2  3  4  CMBH  PARAMS:
+  L1=3.7893m
+  L2=361.3884u
+  L3=33.0498u
+  L4=2.0011u
+  L5=100.2971n
+  C1=14.6694p
+  C2=35.0003p
+  Rs1=27.0621k
+  Rs2=10.0050k
+  Rs3=300.0049
+  Rs4=659.9999
+  Rs5=259.9997
+  R2=1.4100
+  dL3=1.2904u
+  dC3=6.6536p
+  dL4=6.4880n
+  dC4=83.6198p
+  dR3=480.6655m
+  dR4=8.1730k
+  dR5=780.0033m
+  dR6=26.6000k
+  Rdc=37m
+  ck=143f
.ends 
****
.SUBCKT L_744834405_5m  1  2  3  4
X1  1  2  3  4  CMBH  PARAMS:
+  L1=426.7692u
+  L2=496.4710u
+  L3=4.2160m
+  L4=1.0332m
+  L5=299.4135n
+  C1=20.2291p
+  C2=21.4079p
+  Rs1=28.5719k
+  Rs2=2.5909k
+  Rs3=25.8384k
+  Rs4=640.0066k
+  Rs5=236.3219
+  R2=999.9240m
+  dL3=2.1538u
+  dL4=35.8347n
+  dC3=8.5028p
+  dC4=41.0969p
+  dR3=80.0193m
+  dR4=8.8052k
+  dR5=11.0015
+  dR6=9.8509k
+  Rdc=50m
+  ck=385.5f
.ends 
****  
.SUBCKT L_744834407_7m  1  2  3  4
X1  1  2  3  4  CMBH  PARAMS:
+  L1=602.7567u
+  L2=615.5643u
+  L3=5.6145m
+  L4=528.6856u
+  L5=499.7727n
+  C1=15.2392p
+  C2=9.3742p
+  Rs1=2.2694k
+  Rs2=5.5795k
+  Rs3=52.0072k
+  Rs4=540.0004k
+  Rs5=436.3289
+  R2=999.9916m
+  dL3=2.2724u
+  dL4=44.9815n
+  dC3=8.8984p
+  dC4=29.0067p
+  dR3=80.0037m
+  dR4=13.0796k
+  dR5=18.0001
+  dR6=59.8500k
+  Rdc=80m
+  ck=147.8f
.ends  
**** 
.SUBCKT L_744834310_10m  1  2  3  4
X1  1  2  3  4  CMBH  PARAMS:
+  L1=10m
+  L2=250u
+  L3=13u
+  L4=0.1u
+  L5=100.4n
+  C1=12.7p
+  C2=17.2p
+  Rs1=97k
+  Rs2=12k
+  Rs3=200
+  Rs4=260
+  Rs5=460
+  R2=1.41
+  dL3=4.4201u
+  dC3=6.6171p
+  dL4=12.7711n
+  dC4=21.2990p
+  dR3=1.4897
+  dR4=20.0594k
+  dR5=17.0002
+  dR6=866.0004
+  Rdc=110m
+  ck=151.2731f
.ends  
****
.SUBCKT L_744834220_20m  1  2  3  4
X1  1  2  3  4  CMBH  PARAMS:
+  L1=20m
+  L2=250u
+  L3=13u
+  L4=100n
+  L5=100.4n
+  C1=22.2p
+  C2=41.2p
+  Rs1=215k
+  Rs2=2k
+  Rs3=200
+  Rs4=260
+  Rs5=400
+  R2=1.41
+  dL3=7.8522u
+  dC3=11.5456p
+  dL4=652.4980n
+  dC4=162.8939p
+  dR3=489.9657m
+  dR4=27.3787k
+  dR5=1.5000k
+  dR6=8.6600k
+  Rdc=230m
+  ck=103.02f
.ends  
****
.SUBCKT CMBH  1  2  3  4  PARAMS:
R_R9  N12325  3  {R2}
R_R8  N13265  N13287  {Rs4}  
Kn_K6  L_L11  L_L12
+  L_L13  L_L14  0.9999
R_R3  N12571  N12583  {Rs3}
R_R10  N13777  4  {R2}
C_C10  N13029  N12821  {ck}
R_R20  N13215  N13229  {dR4}
L_L11  N12821  N12295  {dL4}
R_R17  N12267  N12273  {dR3}
L_L8  N13265  N13287  {L4}
R_R7  N13287  N13305  {Rs3}
L_L9  N12295  N12307  {L5}
Kn_K4  L_L7  L_L8  1
R_R2  N12583  N12599  {Rs2}
Kn_K5  L_L9  L_L10  1
R_R16  N13229  N13249  {dR6}
Kn_K7  L_L15  L_L16
+  L_L17  L_L18  0.9999
C_C5  N12273  N12289  {dC4}
L_L6  N13287  N13305  {L3}
L_L7  N12307  N12571  {L4}
R_R6  N13305  N13319  {Rs2}
R_R21  1  N12257  {Rdc}
Kn_K3  L_L5  L_L6  1
L_L16  N12257  N12799  {dL3}
C_C8  N13215  N13741  {dC3}
L_L18  N13023  N13215  {dL3}
R_R1  N12599  3  {Rs1}
R_R13  N12289  N12295  {dR5}
L_L4  N13305  N13319  {L2}
L_L5  N12571  N12583  {L3}
R_R15  N13755  N13249  {dR5}
R_R5  N13319  4  {Rs1}
R_R18  N12257  N12273  {dR4}
Kn_K2  L_L3  L_L4  1
R_R19  N13741  N13229  {dR3}
L_L15  N12799  N12273  {dL3}
L_L17  N13229  N13023  {dL3}
L_L3  N12583  N12599  {L2}
R_R11  N12295  N12307  {Rs5}
L_L2  N13319  4  {L1}
C_C4  N13249  N13265  {C2}
L_L10  N13249  N13265  {L5}
Kn_K1  L_L1  L_L2  1
R_R14  N12273  N12295  {dR6}
C_C6  N13229  N13755  {dC4}
L_L12  N12273  N12821  {dL4}
L_L14  N13029  N13229  {dL4}
L_L1  N12599  3  {L1}
C_C1  N12307  N12325  {C1}
R_R12  N13249  N13265  {Rs5}
C_C2  N13265  N13777  {C1}
R_R22  2  N13215  {Rdc}
C_C9  N13023  N12799  {ck}
R_R4  N12307  N12571  {Rs4}
C_C3  N12295  N12307  {C2}
L_L13  N13249  N13029  {dL4}
C_C7  N12257  N12267  {dC3}
.ends  CMBH
****