**************************************************
* Manufacturer:          Würth Elektronik
* Kinds:                 Film Capacitor
* Matchcode:             WCAP-FTDB
* Library Type:          LTspice
* Version:               rev23a
* Created/modified by:   Ella
* Date and Time:         11/22/2023
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2023 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 890764429002CS_60uF 1 2
Rser 1 3 0.0115
Lser 2 4 13.4
C1 3 4 0.00006
Rpar 3 4 166666666.666667
.ends 890764429002CS_60uF
*******
.subckt 890764428004CS_40uF 1 2
Rser 1 3 0.02
Lser 2 4 15.3
C1 3 4 0.00004
Rpar 3 4 250000000
.ends 890764428004CS_40uF
*******
.subckt 890764427009CS_10uF 1 2
Rser 1 3 0.014
Lser 2 4 30
C1 3 4 0.00001
Rpar 3 4 1000000000
.ends 890764427009CS_10uF
*******
.subckt 890744429005CS_40uF 1 2
Rser 1 3 0.017
Lser 2 4 12.2
C1 3 4 0.00004
Rpar 3 4 250000000
.ends 890744429005CS_40uF
*******
.subckt 890744429002CS_25uF 1 2
Rser 1 3 0.021
Lser 2 4 17.3
C1 3 4 0.000025
Rpar 3 4 400000000
.ends 890744429002CS_25uF
*******
.subckt 890744428006CS_25uF 1 2
Rser 1 3 0.0125
Lser 2 4 16.1
C1 3 4 0.000025
Rpar 3 4 400000000
.ends 890744428006CS_25uF
*******
.subckt 890744427005CS_5uF 1 2
Rser 1 3 0.05
Lser 2 4 11.4
C1 3 4 0.000005
Rpar 3 4 2000000000
.ends 890744427005CS_5uF
*******
.subckt 890744427001CS_1uF 1 2
Rser 1 3 0.013
Lser 2 4 13.3
C1 3 4 0.000001
Rpar 3 4 10000000000
.ends 890744427001CS_1uF
*******
.subckt 890734429007CS_50uF 1 2
Rser 1 3 0.0058
Lser 2 4 15.8
C1 3 4 0.00005
Rpar 3 4 200000000
.ends 890734429007CS_50uF
*******
.subckt 890734428008CS_30uF 1 2
Rser 1 3 0.006
Lser 2 4 28.4
C1 3 4 0.00003
Rpar 3 4 333333333.333333
.ends 890734428008CS_30uF
*******
.subckt 890734428004CS_15uF 1 2
Rser 1 3 0.0105
Lser 2 4 32.1
C1 3 4 0.000015
Rpar 3 4 666666666.666667
.ends 890734428004CS_15uF
*******
.subckt 890734427005CS_3uF 1 2
Rser 1 3 0.0075
Lser 2 4 34.9
C1 3 4 0.000003
Rpar 3 4 3333333333.33333
.ends 890734427005CS_3uF
*******
.subckt 890724429010CS_75uF 1 2
Rser 1 3 0.0043
Lser 2 4 41
C1 3 4 0.000075
Rpar 3 4 133333333.333333
.ends 890724429010CS_75uF
*******
.subckt 890724429005CS_50uF 1 2
Rser 1 3 0.007
Lser 2 4 28.7
C1 3 4 0.00005
Rpar 3 4 200000000
.ends 890724429005CS_50uF
*******
.subckt 890724427010CS_10uF 1 2
Rser 1 3 0.016
Lser 2 4 15.5
C1 3 4 0.00001
Rpar 3 4 1000000000
.ends 890724427010CS_10uF
*******
.subckt 890724427001CS_1uF 1 2
Rser 1 3 0.00585153402299
Lser 2 4 25.169149709
C1 3 4 0.000001
Rpar 3 4 10000000000
.ends 890724427001CS_1uF
*******
.subckt 890714429003CS_50uF 1 2
Rser 1 3 0.0082424291924
Lser 2 4 29.391658793
C1 3 4 0.00005
Rpar 3 4 200000000
.ends 890714429003CS_50uF
*******
.subckt 890494429005CS_50uF 1 2
Rser 1 3 0.00613739336009
Lser 2 4 26.31067956
C1 3 4 0.00005
Rpar 3 4 200000000
.ends 890494429005CS_50uF
*******
.subckt 890494429003CS_40uF 1 2
Rser 1 3 0.00693063421548
Lser 2 4 36.302615749
C1 3 4 0.00004
Rpar 3 4 250000000
.ends 890494429003CS_40uF
*******
.subckt 890494428004CS_25uF 1 2
Rser 1 3 0.004
Lser 2 4 32
C1 3 4 0.000025
Rpar 3 4 400000000
.ends 890494428004CS_25uF
*******
.subckt 890494427003CS_3uF 1 2
Rser 1 3 0.00571873831026
Lser 2 4 44.252244217
C1 3 4 0.000003
Rpar 3 4 3333333333.33333
.ends 890494427003CS_3uF
*******
.subckt 890484429001CS_75uF 1 2
Rser 1 3 0.0495
Lser 2 4 13.5
C1 3 4 0.000075
Rpar 3 4 133333333.333333
.ends 890484429001CS_75uF
*******
.subckt 890484428002CS_35uF 1 2
Rser 1 3 0.00654658420506
Lser 2 4 47.8760863
C1 3 4 0.000035
Rpar 3 4 285714285.714286
.ends 890484428002CS_35uF
*******
.subckt 890484427001CS_5uF 1 2
Rser 1 3 0.0047
Lser 2 4 22.8
C1 3 4 0.000005
Rpar 3 4 2000000000
.ends 890484427001CS_5uF
*******
