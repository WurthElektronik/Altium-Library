**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  THT Mono-color Round Color
* Matchcode:              WL-TMRC
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-23
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 3mm_151031SS04000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=1.8860
+ RS=1.0000E-6
+ IKF=1.0000E3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3mm_151031SS06000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=2.0063
+ RS=1.0000E-6
+ IKF=83.795E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3mm_151031VS04000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=1.9467
+ RS=1.0000E-6
+ IKF=16.664E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3mm_151031VS06000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=1.9531
+ RS=1.0000E-6
+ IKF=4.1566E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3mm_151031YS05900  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=1.9096
+ RS=1.0000E-6
+ IKF=5.3812E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3mm_151031YS06000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=1.8193
+ RS=1.0000E-6
+ IKF=16.654E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 5mm_151051BS04000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=2.8744
+ RS=1.0000E-6
+ IKF=4.1539E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 5mm_151051RS11000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=1.9769
+ RS=1.0000E-6
+ IKF=1.0000E3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 5mm_151051SS04000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=1.9451
+ RS=1.0000E-6
+ IKF=1.0000E3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 5mm_151051VS04000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=2.0120
+ RS=1.0000E-6
+ IKF=1.0000E3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 5mm_151051YS04000  1  2
D1 1 2 TMRC
.MODEL TMRC D
+ IS=10.010E-21
+ N=1.9146
+ RS=1.0000E-6
+ IKF=1.0000E3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******






























