**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  Sleeve Choke 
* Matchcode:              WE-WAFB 
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Ella      
* Date and Time:          2022-11-08
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 4535_7427603_70ohm 1 2
Rp 1 2 100
Cp 1 2 0.4p
Rs 1 N3 0.005
L1 N3 2 0.6u
.ends 4535_7427603_70ohm
*******
.subckt 4535_74276031_80ohm 1 2
Rp 1 2 80
Cp 1 2 0.001p
Rs 1 N3 0.005
L1 N3 2 0.42u
.ends 4535_74276031_80ohm
*******
.subckt 5035_74276032_83ohm 1 2
Rp 1 2 105
Cp 1 2 0.2p
Rs 1 N3 0.005
L1 N3 2 0.85u
.ends 5035_74276032_83ohm
*******
.subckt 6035_7427604_82ohm 1 2
Rp 1 2 115
Cp 1 2 0.01p
Rs 1 N3 0.005
L1 N3 2 0.7u
.ends 6035_7427604_82ohm
*******
.subckt 6035_74276041_89ohm 1 2
Rp 1 2 90
Cp 1 2 0.001p
Rs 1 N3 0.005
L1 N3 2 0.72u
.ends 6035_74276041_89ohm
*******
.subckt 7535_7427605_100ohm 1 2
Rp 1 2 135
Cp 1 2 0.05p
Rs 1 N3 0.005
L1 N3 2 0.99u
.ends 7535_7427605_100ohm
*******
.subckt 7835_74276051_100ohm 1 2
Rp 1 2 105
Cp 1 2 0.01p
Rs 1 N3 0.005
L1 N3 2 0.58u
.ends 7835_74276051_100ohm
*******
.subckt 8335_7427602_130ohm 1 2
Rp 1 2 150
Cp 1 2 0.05p
Rs 1 N3 0.005
L1 N3 2 0.85u
.ends 8335_7427602_130ohm
*******
.subckt 9035_7427606_130ohm 1 2
Rp 1 2 130
Cp 1 2 0.01p
Rs 1 N3 0.005
L1 N3 2 1.2u
.ends 9035_7427606_130ohm
*******
.subckt 4535_7427620_130ohm 1 2
Rp 1 2 135
Cp 1 2 0.1p
Rs 1 N3 0.02
L1 N3 2 0.85u
.ends 4535_7427620_130ohm
*******