**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Off-Line Transformer
* Matchcode:              WE-UNIT
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Toby      
* Date and Time:          2022-05-17
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************

.subckt 749118105		3  1  4  6		
.param RxLkg=31788.83ohm					
.param Leakage=150uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	2650uH	Rser=8350mohm	
Lsec1	4	6	7.848uH	Rser=26mohm	
K Lpri1    Lsec1        1					
.param Cprm1=19.88pf					
.param Rdmp1=593391.56ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	1	0	20meg		
Rg11	4	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt 7491181012		3  1  4  6		
.param RxLkg=26640.04ohm					
.param Leakage=134uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	2666uH	Rser=8350mohm	
Lsec1	4	6	42.727uH	Rser=148mohm	
K Lpri1    Lsec1        1					
.param Cprm1=22.59pf					
.param Rdmp1=556657.55ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	1	0	20meg		
Rg11	4	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt 7491181024		3  1  4  6		
.param RxLkg=28569.08ohm					
.param Leakage=145uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	2655uH	Rser=8350mohm	
Lsec1	4	6	170.907uH	Rser=670mohm	
K Lpri1    Lsec1        1					
.param Cprm1=23pf					
.param Rdmp1=551678.75ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	1	0	20meg		
Rg11	4	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt 749118115		5  1  6  9		
.param RxLkg=17392.9ohm					
.param Leakage=87uh					
Rlkg	5	5a	{RxLkg}		
L_Lkg	5	5a	{Leakage}	Rser=0.01mohm	
Lpri1	5a	1	2713uH	Rser=5500mohm	
Lsec1	6	9	7.848uH	Rser=27mohm	
K Lpri1    Lsec1        1					
.param Cprm1=22.34pf					
.param Rdmp1=559771.49ohm					
Cpri1	5	1	{Cprm1}	Rser=10mohm	
Rdmp1	5	1	{Rdmp1}		
Rg3	5	0	20meg		
Rg7	1	0	20meg		
Rg11	6	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt 7491181112		5  1  6  9		
.param RxLkg=16009.14ohm					
.param Leakage=83uh					
Rlkg	5	5a	{RxLkg}		
L_Lkg	5	5a	{Leakage}	Rser=0.01mohm	
Lpri1	5a	1	2717uH	Rser=5500mohm	
Lsec1	6	9	42.727uH	Rser=143mohm	
K Lpri1    Lsec1        1					
.param Cprm1=24pf					
.param Rdmp1=540067.42ohm					
Cpri1	5	1	{Cprm1}	Rser=10mohm	
Rdmp1	5	1	{Rdmp1}		
Rg3	5	0	20meg		
Rg7	1	0	20meg		
Rg11	6	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt 7491181124		5  1  6  9		
.param RxLkg=15788.78ohm					
.param Leakage=81uh					
Rlkg	5	5a	{RxLkg}		
L_Lkg	5	5a	{Leakage}	Rser=0.01mohm	
Lpri1	5a	1	2719uH	Rser=5500mohm	
Lsec1	6	9	170.907uH	Rser=636mohm	
K Lpri1    Lsec1        1					
.param Cprm1=23.5pf					
.param Rdmp1=545785.12ohm					
Cpri1	5	1	{Cprm1}	Rser=10mohm	
Rdmp1	5	1	{Rdmp1}		
Rg3	5	0	20meg		
Rg7	1	0	20meg		
Rg11	6	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt 749118205		8  9  3  4  5  6		
.param RxLkg=45184.55ohm					
.param Leakage=105uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.01mohm	
Lpri1	8a	9	795uH	Rser=3000mohm	
Lsec1	3	4	2.493uH	Rser=21mohm	
Lsec2	5	6	2.493uH	Rser=22mohm	
K Lpri1    Lsec1 Lsec2       1					
.param Cprm1=15pf					
.param Rdmp1=387296.17ohm					
Cpri1	8	9	{Cprm1}	Rser=10mohm	
Rdmp1	8	9	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	9	0	20meg		
Rg11	3	0	20meg		
Rg12	5	0	20meg		
Rg19	4	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt 7491182012		8  9  3  4  5  6		
.param RxLkg=29376.66ohm					
.param Leakage=80uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.01mohm	
Lpri1	8a	9	820uH	Rser=3000mohm	
Lsec1	3	4	9.972uH	Rser=63mohm	
Lsec2	5	6	9.972uH	Rser=70mohm	
K Lpri1    Lsec1 Lsec2       1					
.param Cprm1=20.6pf					
.param Rdmp1=330487.38ohm					
Cpri1	8	9	{Cprm1}	Rser=10mohm	
Rdmp1	8	9	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	9	0	20meg		
Rg11	3	0	20meg		
Rg12	5	0	20meg		
Rg19	4	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt 7491182024		8  9  3  4		
.param RxLkg=28235.13ohm					
.param Leakage=80uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.01mohm	
Lpri1	8a	9	820uH	Rser=3000mohm	
Lsec1	3	4	46.814uH	Rser=180mohm	
K Lpri1    Lsec1        1					
.param Cprm1=22.3pf					
.param Rdmp1=317645.18ohm					
Cpri1	8	9	{Cprm1}	Rser=10mohm	
Rdmp1	8	9	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	9	0	20meg		
Rg11	3	0	20meg		
Rg19	4	0	20meg		
.ends					

.subckt 749118215		3  1  6  7  8  9		
.param RxLkg=20860.31ohm					
.param Leakage=57uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	843uH	Rser=3000mohm	
Lsec1	6	7	2.493uH	Rser=24mohm	
Lsec2	8	9	2.493uH	Rser=25.4mohm	
K Lpri1    Lsec1 Lsec2       1					
.param Cprm1=20.74pf					
.param Rdmp1=329373.37ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	1	0	20meg		
Rg11	6	0	20meg		
Rg12	8	0	20meg		
Rg19	7	0	20meg		
Rg20	9	0	20meg		
.ends					

.subckt 7491182112		3  1  6  7  8  9		
.param RxLkg=18990.39ohm					
.param Leakage=55uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	845uH	Rser=3000mohm	
Lsec1	6	7	9.972uH	Rser=80mohm	
Lsec2	8	9	9.972uH	Rser=87mohm	
K Lpri1    Lsec1 Lsec2       1					
.param Cprm1=23.3pf					
.param Rdmp1=310751.89ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	1	0	20meg		
Rg11	6	0	20meg		
Rg12	8	0	20meg		
Rg19	7	0	20meg		
Rg20	9	0	20meg		
.ends					

.subckt 7491182124		3  1  7  8		
.param RxLkg=17545.17ohm					
.param Leakage=52uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	848uH	Rser=3000mohm	
Lsec1	7	8	46.814uH	Rser=127mohm	
K Lpri1    Lsec1        1					
.param Cprm1=24.4pf					
.param Rdmp1=303666.35ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	1	0	20meg		
Rg11	7	0	20meg		
Rg19	8	0	20meg		
.ends					
