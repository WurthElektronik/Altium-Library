**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT High Current Wire Wound Ceramic Inductor
* Matchcode:              WE-KI HC
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Ella      
* Date and Time:          2022-11-07
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0402_744916010_1n 1 2
C1 1 N7 101.5322f
L1 1 N1 0.95n
L2 N1 N2 64.6465p
L3 N2 N3 86.9525p
L4 N3 N4 28.1671p
L5 N4 N5 62.6356p
L6 N5 N6 49.8196p
R1 2 N1 216.8855m
R2 2 N2 51.4498m
R3 2 N3 47.1552m
R4 2 N4 20.7392m
R5 2 N5 85.3207m
R6 2 N6 68.7325m
R7 2 N7 1.9645
R8 2 1 10g
.ends 
*******
.subckt 0402_744916020_2n 1 2
C1 1 N7 51.2268f
L1 1 N1 1.95n
L2 N1 N2 33.5237p
L3 N2 N3 69.4358p
L4 N3 N4 158.6538p
L5 N4 N5 63.3607p
L6 N5 N6 50.0519p
R1 2 N1 585.5176m
R2 2 N2 324.4036m
R3 2 N3 123.8848m
R4 2 N4 139.6672m
R5 2 N5 85.7777m
R6 2 N6 69.1171m
R7 2 N7 1.965
R8 2 1 10g
.ends 
*******
.subckt 0402_744916022_2.2n 1 2
C1 1 N7 51.5012f
L1 1 N1 2.15n
L2 N1 N2 42.2968p
L3 N2 N3 78.4487p
L4 N3 N4 146.8444p
L5 N4 N5 63.0507p
L6 N5 N6 49.9418p
R1 2 N1 619.9196m
R2 2 N2 367.1853m
R3 2 N3 98.2266m
R4 2 N4 29.4329m
R5 2 N5 84.0186m
R6 2 N6 66.5310m
R7 2 N7 1.9651
R8 2 1 10g
.ends 
*******
.subckt 0402_744916027_2.7n 1 2
C1 1 N7 51.4984f
L1 1 N1 2.6n
L2 N1 N2 42.4697p
L3 N2 N3 94.1194p
L4 N3 N4 153.6619p
L5 N4 N5 63.0625p
L6 N5 N6 49.9456p
R1 2 N1 619.8866m
R2 2 N2 368.9495m
R3 2 N3 105.0213m
R4 2 N4 42.0533m
R5 2 N5 84.0261m
R6 2 N6 66.5377m
R7 2 N7 1.9651
R8 2 1 10g
.ends 
*******
.subckt 0402_744916033_3.3n 1 2
C1 1 N7 53.2352f
L1 1 N1 3.2n
L2 N1 N2 59.9023p
L3 N2 N3 115.2769p
L4 N3 N4 199.9013p
L5 N4 N5 63.2349p
L6 N5 N6 50.0149p
R1 2 N1 724.5164m
R2 2 N2 422.1312m
R3 2 N3 132.3077m
R4 2 N4 118.5406m
R5 2 N5 84.2488m
R6 2 N6 66.8135m
R7 2 N7 1.9657
R8 2 1 10g
.ends 
*******
.subckt 0402_744916036_3.6n 1 2
C1 1 N7 57.5514f
L1 1 N1 3.5n
L2 N1 N2 85.6628p
L3 N2 N3 145.7193p
L4 N3 N4 643.4729p
L5 N4 N5 66.7691p
L6 N5 N6 51.2738p
R1 2 N1 767.5341m
R2 2 N2 538.0661m
R3 2 N3 224.7437m
R4 2 N4 347.1280m
R5 2 N5 96.0084m
R6 2 N6 82.7576m
R7 2 N7 1.9674
R8 2 1 10g
.ends 
*******
.subckt 0402_744916039_3.9n 1 2
C1 1 N7 71.7689f
L1 1 N1 3.8n
L2 N1 N2 86.2701p
L3 N2 N3 108.2969p
L4 N3 N4 642.3604p
L5 N4 N5 66.7612p
L6 N5 N6 51.2715p
R1 2 N1 782.6244m
R2 2 N2 535.8630m
R3 2 N3 212.4643m
R4 2 N4 346.6377m
R5 2 N5 95.9483m
R6 2 N6 82.6798m
R7 2 N7 1.9674
R8 2 1 10g
.ends 
*******
.subckt 0402_744916043_4.3n 1 2
C1 1 N7 97.4069f
L1 1 N1 4.2n
L2 N1 N2 84.1368p
L3 N2 N3 102.8191p
L4 N3 N4 639.1551p
L5 N4 N5 66.7362p
L6 N5 N6 51.2618p
R1 2 N1 750.6952m
R2 2 N2 520.1059m
R3 2 N3 200.9189m
R4 2 N4 346.6254m
R5 2 N5 95.9764m
R6 2 N6 82.7242m
R7 2 N7 1.9673
R8 2 1 10g
.ends 
*******
.subckt 0402_744916047_4.7n 1 2
C1 1 N7 114.8f
L1 1 N1 4.6n
L2 N1 N2 13.3244p
L3 N2 N3 67.8420p
L4 N3 N4 176.8400p
L5 N4 N5 77.3771p
L6 N5 N6 55.1411p
R1 2 N1 2.4046
R2 2 N2 1.2078
R3 2 N3 913.5711m
R4 2 N4 731.8989m
R5 2 N5 603.2267m
R6 2 N6 592.1230m
R7 2 N7 2.0856
R8 2 1 10g
.ends 
*******
.subckt 0402_744916051_5.1n 1 2
C1 1 N7 107.4f
L1 1 N1 5n
L2 N1 N2 13.3836p
L3 N2 N3 62.0266p
L4 N3 N4 282.7699p
L5 N4 N5 77.4303p
L6 N5 N6 55.1482p
R1 2 N1 2.804
R2 2 N2 2.0053
R3 2 N3 909.4285m
R4 2 N4 733.4708m
R5 2 N5 605.0706m
R6 2 N6 593.7937m
R7 2 N7 2.8865
R8 2 1 10g
.ends 
*******
.subckt 0402_744916056_5.6n 1 2
C1 1 N7 134.1332f
L1 1 N1 5.48n
L2 N1 N2 18.4075p
L3 N2 N3 192.2062p
L4 N3 N4 431.2415p
L5 N4 N5 169.8016p
L6 N5 N6 139.7105p
R1 2 N1 2.4420
R2 2 N2 987.9505m
R3 2 N3 250.0718m
R4 2 N4 81.5229m
R5 2 N5 412.8570m
R6 2 N6 59.5957m
R7 2 N7 2.9100
R8 2 1 10g
.ends 
*******
.subckt 0402_744916062_6.2n 1 2
C1 1 N7 125.2609f
L1 1 N1 6n
L2 N1 N2 132.0124p
L3 N2 N3 141.1686p
L4 N3 N4 914.7352p
L5 N4 N5 85.5011p
L6 N5 N6 58.5019p
R1 2 N1 1.0297
R2 2 N2 1.1604
R3 2 N3 398.1095m
R4 2 N4 598.0355m
R5 2 N5 137.8175m
R6 2 N6 130.5588m
R7 2 N7 1.9588
R8 2 1 10g
.ends 
*******
.subckt 0402_744916068_6.8n 1 2
C1 1 N7 110.0945f
L1 1 N1 6.6n
L2 N1 N2 131.7166p
L3 N2 N3 141.4732p
L4 N3 N4 891.1165p
L5 N4 N5 85.3315p
L6 N5 N6 58.4672p
R1 2 N1 1.0182
R2 2 N2 1.1584
R3 2 N3 333.1323m
R4 2 N4 596.3063m
R5 2 N5 137.6346m
R6 2 N6 130.3905m
R7 2 N7 1.9585
R8 2 1 10g
.ends 
*******
.subckt 0402_744916082_8.2n 1 2
C1 1 N7 129.7857f
L1 1 N1 8n
L2 N1 N2 131.5767p
L3 N2 N3 197.9265p
L4 N3 N4 862.4179p
L5 N4 N5 86.2118p
L6 N5 N6 59.3493p
R1 2 N1 1.6809
R2 2 N2 1.6431
R3 2 N3 499.4604m
R4 2 N4 655.7044m
R5 2 N5 149.7811m
R6 2 N6 143.4479m
R7 2 N7 1.9562
R8 2 1 10g
.ends 
*******
.subckt 0402_744916087_8.7n 1 2
C1 1 N7 111.5704f
L1 1 N1 8.45n
L2 N1 N2 132.9522p
L3 N2 N3 266.6644p
L4 N3 N4 1.5800n
L5 N4 N5 92.9958p
L6 N5 N6 61.5468p
R1 2 N1 1.584
R2 2 N2 2.1555
R3 2 N3 546.4118m
R4 2 N4 860.1517m
R5 2 N5 188.6401m
R6 2 N6 183.6925m
R7 2 N7 1.967
R8 2 1 10g
.ends 
*******
.subckt 0402_744916090_9n 1 2
C1 1 N7 111.5546f
L1 1 N1 8.75n
L2 N1 N2 131.5726p
L3 N2 N3 264.0921p
L4 N3 N4 1.5520n
L5 N4 N5 92.7896p
L6 N5 N6 61.5016p
R1 2 N1 1.5001
R2 2 N2 2.1225
R3 2 N3 369.4164m
R4 2 N4 859.1265m
R5 2 N5 188.5583m
R6 2 N6 183.6387m
R7 2 N7 1.9684
R8 2 1 10g
.ends 
*******
.subckt 0402_744916095_9.5n 1 2
C1 1 N7 136.8830f
L1 1 N1 9.25n
L2 N1 N2 131.5734p
L3 N2 N3 289.5965p
L4 N3 N4 1.6134n
L5 N4 N5 93.4838p
L6 N5 N6 61.8791p
R1 2 N1 1.9668
R2 2 N2 2.3534
R3 2 N3 607.8814m
R4 2 N4 884.5296m
R5 2 N5 193.4520m
R6 2 N6 188.6858m
R7 2 N7 1.9655
R8 2 1 10g
.ends 
*******
.subckt 0402_744916110_10n 1 2
C1 1 N7 122.0915f
L1 1 N1 9.7n
L2 N1 N2 131.3909p
L3 N2 N3 289.1961p
L4 N3 N4 1.5966n
L5 N4 N5 93.3703p
L6 N5 N6 61.8596p
R1 2 N1 1.9435
R2 2 N2 2.3418
R3 2 N3 510.0368m
R4 2 N4 885.6048m
R5 2 N5 193.7621m
R6 2 N6 189.0279m
R7 2 N7 1.9662
R8 2 1 10g
.ends 
*******
.subckt 0402_744916111_11n 1 2
C1 1 N7 118.1426f
L1 1 N1 10.65n
L2 N1 N2 120.0986p
L3 N2 N3 321.5246p
L4 N3 N4 1.3227n
L5 N4 N5 91.2436p
L6 N5 N6 61.3813p
R1 2 N1 2.2019
R2 2 N2 2.5381
R3 2 N3 476.0532m
R4 2 N4 870.3854m
R5 2 N5 191.7849m
R6 2 N6 187.2829m
R7 2 N7 1.9672
R8 2 1 10g
.ends 
*******
.subckt 0402_744916112_12n 1 2
C1 1 N7 116.4237f
L1 1 N1 11.65n
L2 N1 N2 19.5700p
L3 N2 N3 510.8978p
L4 N3 N4 3.1352n
L5 N4 N5 99.9596p
L6 N5 N6 64.1561p
R1 2 N1 3.3619
R2 2 N2 2.5503
R3 2 N3 820.8924m
R4 2 N4 1.1158
R5 2 N5 367.7207m
R6 2 N6 365.9667m
R7 2 N7 2.976
R8 2 1 10g
.ends 
*******
.subckt 0402_744916113_13n 1 2
C1 1 N7 126.8346f
L1 1 N1 12.65n
L2 N1 N2 153.8132p
L3 N2 N3 578.7503p
L4 N3 N4 3.0277n
L5 N4 N5 99.9529p
L6 N5 N6 64.1548p
R1 2 N1 3.3723
R2 2 N2 2.5687
R3 2 N3 811.9928m
R4 2 N4 1.1162
R5 2 N5 371.4514m
R6 2 N6 369.7857m
R7 2 N7 2.976
R8 2 1 10g
.ends 
*******
.subckt 0402_744916115_15n 1 2
C1 1 N7 103.2394f
L1 1 N1 14.6n
L2 N1 N2 282.3218p
L3 N2 N3 525.5003p
L4 N3 N4 1.2916n
L5 N4 N5 99.8270p
L6 N5 N6 64.1170p
R1 2 N1 3.382
R2 2 N2 2.5777
R3 2 N3 698.5812m
R4 2 N4 1.1142
R5 2 N5 357.6777m
R6 2 N6 356.9007m
R7 2 N7 2.976
R8 2 1 10g
.ends 
*******
.subckt 0402_744916116_16n 1 2
C1 1 N7 108.0120f
L1 1 N1 15.55n
L2 N1 N2 326.1256p
L3 N2 N3 626.4780p
L4 N3 N4 3.3470n
L5 N4 N5 99.9736p
L6 N5 N6 64.1508p
R1 2 N1 3.3778
R2 2 N2 2.585
R3 2 N3 775.9664m
R4 2 N4 1.1192
R5 2 N5 398.9255m
R6 2 N6 397.1570m
R7 2 N7 2.9762
R8 2 1 10g
.ends 
*******
.subckt 0402_744916118_18n 1 2
C1 1 N7 108.2189f
L1 1 N1 17.55n
L2 N1 N2 388.2772p
L3 N2 N3 635.1311p
L4 N3 N4 3.0901n
L5 N4 N5 99.9555p
L6 N5 N6 64.1464p
R1 2 N1 3.3835
R2 2 N2 2.5907
R3 2 N3 763.9195m
R4 2 N4 1.119
R5 2 N5 397.3205m
R6 2 N6 395.6814m
R7 2 N7 2.9763
R8 2 1 10g
.ends 
*******
.subckt 0402_744916119_19n 1 2
C1 1 N7 100.6697f
L1 1 N1 18.55n
L2 N1 N2 466.1262p
L3 N2 N3 709.6348p
L4 N3 N4 3.0124n
L5 N4 N5 89.3353p
L6 N5 N6 64.1598p
R1 2 N1 4.313
R2 2 N2 2.5331
R3 2 N3 1.7409
R4 2 N4 2.1427
R5 2 N5 681.4697m
R6 2 N6 680.7511m
R7 2 N7 3.2661
R8 2 1 10g
.ends 
*******
.subckt 0402_744916121_21n 1 2
C1 1 N7 101.8489f
L1 1 N1 20.5n
L2 N1 N2 588.4391p
L3 N2 N3 730.8236p
L4 N3 N4 2.6789n
L5 N4 N5 87.7404p
L6 N5 N6 64.1623p
R1 2 N1 4.3157
R2 2 N2 2.549
R3 2 N3 1.728
R4 2 N4 2.1444
R5 2 N5 698.1719m
R6 2 N6 697.5749m
R7 2 N7 3.2653
R8 2 1 10g
.ends 
*******
.subckt 0402_744916122_22n 1 2
C1 1 N7 91.3860f
L1 1 N1 21.2n
L2 N1 N2 515.9474p
L3 N2 N3 768.2286p
L4 N3 N4 3.7453n
L5 N4 N5 96.3660p
L6 N5 N6 64.1863p
R1 2 N1 4.2774
R2 2 N2 3.5618
R3 2 N3 1.7241
R4 2 N4 2.1492
R5 2 N5 740.6104m
R6 2 N6 739.7216m
R7 2 N7 4.2614
R8 2 1 10g
.ends 
*******
.subckt 0402_744916123_23n 1 2
C1 1 N7 100.1717f
L1 1 N1 22.2n
L2 N1 N2 719.0542p
L3 N2 N3 904.2044p
L4 N3 N4 5.7324n
L5 N4 N5 105.2278p
L6 N5 N6 64.2049p
R1 2 N1 3.5913
R2 2 N2 2.6452
R3 2 N3 1.0068
R4 2 N4 1.1361
R5 2 N5 505.1302m
R6 2 N6 503.0742m
R7 2 N7 4.2778
R8 2 1 10g
.ends 
*******
.subckt 0402_744916124_24n 1 2
C1 1 N7 104.7791f
L1 1 N1 23.2n
L2 N1 N2 881.7684p
L3 N2 N3 913.2233p
L4 N3 N4 5.6069n
L5 N4 N5 106.2006p
L6 N5 N6 64.2325p
R1 2 N1 3.6315
R2 2 N2 2.6592
R3 2 N3 998.4371m
R4 2 N4 1.1372
R5 2 N5 510.4903m
R6 2 N6 508.5292m
R7 2 N7 4.2789
R8 2 1 10g
.ends 
*******
.subckt 0402_744916125_25n 1 2
C1 1 N7 99.0782f
L1 1 N1 24.2n
L2 N1 N2 881.7272p
L3 N2 N3 913.1728p
L4 N3 N4 5.6061n
L5 N4 N5 106.2057p
L6 N5 N6 64.2327p
R1 2 N1 3.6315
R2 2 N2 2.6592
R3 2 N3 998.3715m
R4 2 N4 1.1372
R5 2 N5 510.5229m
R6 2 N6 508.5624m
R7 2 N7 4.2789
R8 2 1 10g
.ends 
*******
.subckt 0402_744916126_26n 1 2
C1 1 N7 91.9644f
L1 1 N1 25.1n
L2 N1 N2 658.6573p
L3 N2 N3 795.3333p
L4 N3 N4 3.6339n
L5 N4 N5 96.1355p
L6 N5 N6 64.1926p
R1 2 N1 4.2947
R2 2 N2 3.5746
R3 2 N3 1.7218
R4 2 N4 2.1494
R5 2 N5 742.2699m
R6 2 N6 741.4173m
R7 2 N7 4.2627
R8 2 1 10g
.ends 
*******
.subckt 0402_744916127_27n 1 2
C1 1 N7 88.3320f
L1 1 N1 26.1n
L2 N1 N2 681.8502p
L3 N2 N3 762.7428p
L4 N3 N4 2.6714n
L5 N4 N5 89.9138p
L6 N5 N6 64.1806p
R1 2 N1 4.2966
R2 2 N2 3.5707
R3 2 N3 1.684
R4 2 N4 2.1511
R5 2 N5 757.4297m
R6 2 N6 756.8736m
R7 2 N7 4.2623
R8 2 1 10g
.ends 
*******
.subckt 0402_744916130_30n 1 2
C1 1 N7 77.5919f
L1 1 N1 29n
L2 N1 N2 1.0587n
L3 N2 N3 687.8073p
L4 N3 N4 3.4363n
L5 N4 N5 98.1794p
L6 N5 N6 64.2192p
R1 2 N1 4.4806
R2 2 N2 3.5774
R3 2 N3 1.6454
R4 2 N4 2.1609
R5 2 N5 830.0149m
R6 2 N6 829.2924m
R7 2 N7 4.2813
R8 2 1 10g
.ends 
*******
.subckt 0402_744916133_33n 1 2
C1 1 N7 76.9569f
L1 1 N1 32n
L2 N1 N2 1.1638n
L3 N2 N3 672.6417p
L4 N3 N4 6.8640n
L5 N4 N5 125.7485p
L6 N5 N6 64.3285p
R1 2 N1 5.3476
R2 2 N2 3.603
R3 2 N3 2.039
R4 2 N4 2.2339
R5 2 N5 1.2318
R6 2 N6 1.2312
R7 2 N7 4.4201
R8 2 1 10g
.ends 
*******
.subckt 0402_744916136_36n 1 2
C1 1 N7 77.1246f
L1 1 N1 34.9n
L2 N1 N2 1.2321n
L3 N2 N3 663.3121p
L4 N3 N4 4.4423n
L5 N4 N5 111.2809p
L6 N5 N6 64.2988p
R1 2 N1 5.3667
R2 2 N2 3.5913
R3 2 N3 1.9801
R4 2 N4 2.2325
R5 2 N5 1.2288
R6 2 N6 1.2286
R7 2 N7 4.4242
R8 2 1 10g
.ends 
*******
.subckt 0402_744916137_37n 1 2
C1 1 N7 68.6866f
L1 1 N1 35.9n
L2 N1 N2 1.4891n
L3 N2 N3 644.9443p
L4 N3 N4 4.9391n
L5 N4 N5 116.4861p
L6 N5 N6 64.3351p
R1 2 N1 5.6857
R2 2 N2 3.8118
R3 2 N3 2.2421
R4 2 N4 2.2693
R5 2 N5 1.3422
R6 2 N6 1.342
R7 2 N7 4.4705
R8 2 1 10g
.ends 
*******
.subckt 0402_744916139_39n 1 2
C1 1 N7 64.8819f
L1 1 N1 37.7n
L2 N1 N2 1.4780n
L3 N2 N3 618.1339p
L4 N3 N4 5.0570n
L5 N4 N5 102.3034p
L6 N5 N6 64.1699p
R1 2 N1 5.5438
R2 2 N2 3.4878
R3 2 N3 3.8416
R4 2 N4 2.1839
R5 2 N5 900.5737m
R6 2 N6 899.8789m
R7 2 N7 7.9599
R8 2 1 10g
.ends 
*******
.subckt 0402_744916140_40n 1 2
C1 1 N7 70.2538f
L1 1 N1 38.5n
L2 N1 N2 1.0484n
L3 N2 N3 964.4523p
L4 N3 N4 2.5743n
L5 N4 N5 69.5174p
L6 N5 N6 63.6368p
R1 2 N1 7.9537
R2 2 N2 4.0171
R3 2 N3 4.3263
R4 2 N4 2.6803
R5 2 N5 2.1552
R6 2 N6 2.1554
R7 2 N7 9.2825
R8 2 1 10g
.ends 
*******
.subckt 0402_744916143_43n 1 2
C1 1 N7 60.8640f
L1 1 N1 41.5n
L2 N1 N2 1.4824n
L3 N2 N3 366.7905p
L4 N3 N4 3.6044n
L5 N4 N5 75.2082p
L6 N5 N6 63.6374p
R1 2 N1 8.2671
R2 2 N2 3.744
R3 2 N3 4.128
R4 2 N4 2.6796
R5 2 N5 2.1543
R6 2 N6 2.1543
R7 2 N7 9.3704
R8 2 1 10g
.ends 
*******
.subckt 0402_744916147_47n 1 2
C1 1 N7 65.2771f
L1 1 N1 45.5n
L2 N1 N2 1.6780n
L3 N2 N3 349.8298p
L4 N3 N4 5.1723n
L5 N4 N5 81.4176p
L6 N5 N6 63.6316p
R1 2 N1 8.3405
R2 2 N2 3.7352
R3 2 N3 4.1166
R4 2 N4 2.6838
R5 2 N5 2.1605
R6 2 N6 2.1604
R7 2 N7 9.3829
R8 2 1 10g
.ends 
*******
.subckt 0402_744916151_51n 1 2
C1 1 N7 61.9055f
L1 1 N1 49.5n
L2 N1 N2 2.3730n
L3 N2 N3 323.4464p
L4 N3 N4 6.0706n
L5 N4 N5 106.0228p
L6 N5 N6 63.9856p
R1 2 N1 8.2311
R2 2 N2 3.5013
R3 2 N3 3.8993
R4 2 N4 2.5328
R5 2 N5 1.9081
R6 2 N6 1.9079
R7 2 N7 9.3016
R8 2 1 10g
.ends 
*******
.subckt 0603_744917018_1.8n 1 2
C1 1 N7 50.2250f
L1 1 N1 1.75n
L2 N1 N2 49.0712p
L3 N2 N3 75.5513p
L4 N3 N4 137.5197p
L5 N4 N5 63.3637p
L6 N5 N6 50.0987p
R1 2 N1 621.9681m
R2 2 N2 466.3613m
R3 2 N3 180.9765m
R4 2 N4 139.0182m
R5 2 N5 85.9155m
R6 2 N6 69.3047m
R7 2 N7 1.9651
R8 2 1 10g
.ends 
*******
.subckt 0603_744917022_2.2n 1 2
C1 1 N7 51.1233f
L1 1 N1 2n
L2 N1 N2 87.6443p
L3 N2 N3 125.4170p
L4 N3 N4 816.7157p
L5 N4 N5 70.8219p
L6 N5 N6 53.1271p
R1 2 N1 910.0419m
R2 2 N2 456.8994m
R3 2 N3 93.9877m
R4 2 N4 518.6485m
R5 2 N5 213.1334m
R6 2 N6 209.0448m
R7 2 N7 3.5676
R8 2 1 10g
.ends 
*******
.subckt 0603_744917033_3.3n 1 2
C1 1 N7 46.8538f
L1 1 N1 3.2n
L2 N1 N2 59.2647p
L3 N2 N3 266.0834p
L4 N3 N4 819.1104p
L5 N4 N5 70.7902p
L6 N5 N6 53.0692p
R1 2 N1 660.8300m
R2 2 N2 325.5016m
R3 2 N3 97.5625m
R4 2 N4 518.1386m
R5 2 N5 211.4953m
R6 2 N6 207.2315m
R7 2 N7 3.5667
R8 2 1 10g
.ends 
*******
.subckt 0603_744917036_3.6n 1 2
C1 1 N7 48.6210f
L1 1 N1 3.55n
L2 N1 N2 67.9022p
L3 N2 N3 201.3157p
L4 N3 N4 819.0550p
L5 N4 N5 70.8003p
L6 N5 N6 53.0836p
R1 2 N1 743.3446m
R2 2 N2 340.5208m
R3 2 N3 97.3400m
R4 2 N4 518.1794m
R5 2 N5 211.2383m
R6 2 N6 206.9667m
R7 2 N7 3.5672
R8 2 1 10g
.ends 
*******
.subckt 0603_744917039_3.9n 1 2
C1 1 N7 52.8754f
L1 1 N1 3.8n
L2 N1 N2 83.3504p
L3 N2 N3 191.8094p
L4 N3 N4 793.4875p
L5 N4 N5 70.6308p
L6 N5 N6 53.0524p
R1 2 N1 891.1123m
R2 2 N2 377.6745m
R3 2 N3 92.5677m
R4 2 N4 513.3461m
R5 2 N5 186.0691m
R6 2 N6 183.2017m
R7 2 N7 3.5683
R8 2 1 10g
.ends 
*******
.subckt 0603_744917043_4.3n 1 2
C1 1 N7 60.4785f
L1 1 N1 4.2n
L2 N1 N2 108.0239p
L3 N2 N3 232.5395p
L4 N3 N4 685.0326p
L5 N4 N5 69.8378p
L6 N5 N6 52.8728p
R1 2 N1 1.0981
R2 2 N2 432.5323m
R3 2 N3 76.9517m
R4 2 N4 498.0933m
R5 2 N5 77.9540m
R6 2 N6 86.3507m
R7 2 N7 3.5704
R8 2 1 10g
.ends 
*******
.subckt 0603_744917051_5.1n 1 2
C1 1 N7 47.9035f
L1 1 N1 5n
L2 N1 N2 98.9541p
L3 N2 N3 302.3313p
L4 N3 N4 831.8527p
L5 N4 N5 70.9066p
L6 N5 N6 53.1352p
R1 2 N1 893.0466m
R2 2 N2 500.1877m
R3 2 N3 113.4822m
R4 2 N4 515.6299m
R5 2 N5 228.3377m
R6 2 N6 218.2817m
R7 2 N7 3.5661
R8 2 1 10g
.ends 
*******
.subckt 0603_744917056_5.6n 1 2
C1 1 N7 103.3733f
L1 1 N1 5.45n
L2 N1 N2 115.1884p
L3 N2 N3 215.0997p
L4 N3 N4 758.0070p
L5 N4 N5 70.3644p
L6 N5 N6 53.0033p
R1 2 N1 875.5592m
R2 2 N2 462.2488m
R3 2 N3 105.4456m
R4 2 N4 498.2630m
R5 2 N5 88.3103m
R6 2 N6 39.9342m
R7 2 N7 1.5725
R8 2 1 10g
.ends 
*******
.subckt 0603_744917060_6n 1 2
C1 1 N7 118.8660f
L1 1 N1 5.85n
L2 N1 N2 99.9318p
L3 N2 N3 309.3061p
L4 N3 N4 812.8811p
L5 N4 N5 70.7974p
L6 N5 N6 53.1230p
R1 2 N1 1.0448
R2 2 N2 417.4356m
R3 2 N3 114.3534m
R4 2 N4 504.4716m
R5 2 N5 167.5605m
R6 2 N6 174.9210m
R7 2 N7 1.5844
R8 2 1 10g
.ends 
*******
.subckt 0603_744917068_6.8n 1 2
C1 1 N7 110.9262f
L1 1 N1 6.6n
L2 N1 N2 119.7323p
L3 N2 N3 430.5137p
L4 N3 N4 861.4979p
L5 N4 N5 71.1492p
L6 N5 N6 53.2244p
R1 2 N1 1.2224
R2 2 N2 456.7872m
R3 2 N3 124.2220m
R4 2 N4 511.4972m
R5 2 N5 205.9332m
R6 2 N6 206.9738m
R7 2 N7 1.5957
R8 2 1 10g
.ends 
*******
.subckt 0603_744917072_7.2n 1 2
C1 1 N7 120.8179f
L1 1 N1 7n
L2 N1 N2 127.7025p
L3 N2 N3 347.0444p
L4 N3 N4 857.2987p
L5 N4 N5 71.0840p
L6 N5 N6 53.2015p
R1 2 N1 1.233
R2 2 N2 474.7079m
R3 2 N3 128.0162m
R4 2 N4 398.2920m
R5 2 N5 97.2904m
R6 2 N6 91.4828m
R7 2 N7 1.1597
R8 2 1 10g
.ends 
*******
.subckt 0603_744917075_7.5n 1 2
C1 1 N7 126.0059f
L1 1 N1 7.3n
L2 N1 N2 139.9131p
L3 N2 N3 341.4159p
L4 N3 N4 880.9203p
L5 N4 N5 71.2804p
L6 N5 N6 53.2748p
R1 2 N1 1.3072
R2 2 N2 579.6861m
R3 2 N3 131.1534m
R4 2 N4 404.5181m
R5 2 N5 156.4148m
R6 2 N6 152.0720m
R7 2 N7 1.606
R8 2 1 10g
.ends 
*******
.subckt 0603_744917082_8.2n 1 2
C1 1 N7 88.8273f
L1 1 N1 8n
L2 N1 N2 127.6302p
L3 N2 N3 434.7847p
L4 N3 N4 1.2476n
L5 N4 N5 73.4297p
L6 N5 N6 53.8739p
R1 2 N1 1.1298
R2 2 N2 716.8081m
R3 2 N3 189.9458m
R4 2 N4 525.8908m
R5 2 N5 431.5948m
R6 2 N6 420.7209m
R7 2 N7 1.5992
R8 2 1 10g
.ends 
*******
.subckt 0603_744917087_8.7n 1 2
C1 1 N7 92.2899f
L1 1 N1 8.5n
L2 N1 N2 137.5760p
L3 N2 N3 327.1900p
L4 N3 N4 1.2092n
L5 N4 N5 73.2572p
L6 N5 N6 53.8106p
R1 2 N1 1.081
R2 2 N2 482.0759m
R3 2 N3 184.4874m
R4 2 N4 278.8427m
R5 2 N5 399.9369m
R6 2 N6 388.3470m
R7 2 N7 1.1725
R8 2 1 10g
.ends 
*******
.subckt 0603_744917091_9.1n 1 2
C1 1 N7 101.8144f
L1 1 N1 8.9n
L2 N1 N2 159.4457p
L3 N2 N3 731.0274p
L4 N3 N4 1.7925n
L5 N4 N5 75.8757p
L6 N5 N6 54.7351p
R1 2 N1 1.4766
R2 2 N2 809.5875m
R3 2 N3 376.6998m
R4 2 N4 720.8410m
R5 2 N5 716.7037m
R6 2 N6 706.0716m
R7 2 N7 3.4854
R8 2 1 10g
.ends 
*******
.subckt 0603_744917095_9.5n 1 2
C1 1 N7 154.8037f
L1 1 N1 9.3n
L2 N1 N2 158.7972p
L3 N2 N3 294.6232p
L4 N3 N4 956.7403p
L5 N4 N5 72.8164p
L6 N5 N6 53.8485p
R1 2 N1 1.1673
R2 2 N2 505.9899m
R3 2 N3 306.5498m
R4 2 N4 51.4901m
R5 2 N5 134.3688m
R6 2 N6 110.2504m
R7 2 N7 1.6001
R8 2 1 10g
.ends 
*******
.subckt 0603_744917110_10n 1 2
C1 1 N7 174.4643f
L1 1 N1 9.7n
L2 N1 N2 178.5665p
L3 N2 N3 293.8993p
L4 N3 N4 954.5733p
L5 N4 N5 72.8238p
L6 N5 N6 53.8503p
R1 2 N1 1.4123
R2 2 N2 671.6701m
R3 2 N3 305.9432m
R4 2 N4 126.9830m
R5 2 N5 150.0716m
R6 2 N6 132.3369m
R7 2 N7 1.6361
R8 2 1 10g
.ends 
*******
.subckt 0603_744917111_11n 1 2
C1 1 N7 138.5036f
L1 1 N1 10.6n
L2 N1 N2 218.8170p
L3 N2 N3 526.1060p
L4 N3 N4 1.2865n
L5 N4 N5 74.4133p
L6 N5 N6 54.3551p
R1 2 N1 1.7654
R2 2 N2 952.5632m
R3 2 N3 318.0323m
R4 2 N4 481.3113m
R5 2 N5 461.8282m
R6 2 N6 454.3676m
R7 2 N7 1.5909
R8 2 1 10g
.ends 
*******
.subckt 0603_744917112_12n 1 2
C1 1 N7 138.0255f
L1 1 N1 11.6n
L2 N1 N2 235.7715p
L3 N2 N3 680.7955p
L4 N3 N4 1.4206n
L5 N4 N5 75.0490p
L6 N5 N6 54.5530p
R1 2 N1 1.9738
R2 2 N2 921.9259m
R3 2 N3 328.2626m
R4 2 N4 552.8259m
R5 2 N5 530.2108m
R6 2 N6 521.6200m
R7 2 N7 3.6138
R8 2 1 10g
.ends 
*******
.subckt 0603_744917115_15n 1 2
C1 1 N7 130.7211f
L1 1 N1 14.5n
L2 N1 N2 254.1467p
L3 N2 N3 552.0317p
L4 N3 N4 1.4270n
L5 N4 N5 75.1438p
L6 N5 N6 54.6495p
R1 2 N1 2.1205
R2 2 N2 1.1393
R3 2 N3 327.9050m
R4 2 N4 545.5872m
R5 2 N5 521.8682m
R6 2 N6 512.8175m
R7 2 N7 3.6115
R8 2 1 10g
.ends 
*******
.subckt 0603_744917116_16n 1 2
C1 1 N7 128.3145f
L1 1 N1 15.5n
L2 N1 N2 271.7300p
L3 N2 N3 482.3228p
L4 N3 N4 1.2627n
L5 N4 N5 74.3262p
L6 N5 N6 54.4195p
R1 2 N1 2.301
R2 2 N2 1.1982
R3 2 N3 320.2854m
R4 2 N4 238.1587m
R5 2 N5 160.5766m
R6 2 N6 123.4352m
R7 2 N7 3.6214
R8 2 1 10g
.ends 
*******
.subckt 0603_744917118_18n 1 2
C1 1 N7 120.5990f
L1 1 N1 17.5n
L2 N1 N2 359.7126p
L3 N2 N3 1.1079n
L4 N3 N4 2.1411n
L5 N4 N5 78.3308p
L6 N5 N6 55.4300p
R1 2 N1 3.0141
R2 2 N2 1.0028
R3 2 N3 377.2476m
R4 2 N4 925.9245m
R5 2 N5 887.5947m
R6 2 N6 852.3160m
R7 2 N7 3.7099
R8 2 1 10g
.ends 
*******
.subckt 0603_744917122_22n 1 2
C1 1 N7 119.1066f
L1 1 N1 21.5n
L2 N1 N2 438.5944p
L3 N2 N3 1.0768n
L4 N3 N4 2.3040n
L5 N4 N5 79.2270p
L6 N5 N6 55.8381p
R1 2 N1 3.6072
R2 2 N2 1.2174
R3 2 N3 400.9837m
R4 2 N4 912.4685m
R5 2 N5 866.1335m
R6 2 N6 826.3448m
R7 2 N7 3.8341
R8 2 1 10g
.ends 
*******
.subckt 0603_744917123_23n 1 2
C1 1 N7 112.2262f
L1 1 N1 22.4n
L2 N1 N2 538.6750p
L3 N2 N3 1.2184n
L4 N3 N4 2.5378n
L5 N4 N5 80.2989p
L6 N5 N6 56.1105p
R1 2 N1 4.3746
R2 2 N2 1.2574
R3 2 N3 437.2993m
R4 2 N4 882.1871m
R5 2 N5 822.3233m
R6 2 N6 774.1846m
R7 2 N7 4.0431
R8 2 1 10g
.ends 
*******
.subckt 0603_744917124_24n 1 2
C1 1 N7 121.3205f
L1 1 N1 23.4n
L2 N1 N2 429.1656p
L3 N2 N3 884.3258p
L4 N3 N4 2.2055n
L5 N4 N5 78.5969p
L6 N5 N6 55.5475p
R1 2 N1 4.345
R2 2 N2 1.1296
R3 2 N3 394.8550m
R4 2 N4 435.3389m
R5 2 N5 274.9415m
R6 2 N6 133.8933m
R7 2 N7 4.0811
R8 2 1 10g
.ends 
*******
.subckt 0603_744917127_27n 1 2
C1 1 N7 108.0772f
L1 1 N1 26.4n
L2 N1 N2 528.5768p
L3 N2 N3 1.2921n
L4 N3 N4 2.7477n
L5 N4 N5 81.5983p
L6 N5 N6 56.6513p
R1 2 N1 4.7523
R2 2 N2 1.3374
R3 2 N3 447.5840m
R4 2 N4 723.0013m
R5 2 N5 808.6818m
R6 2 N6 771.7510m
R7 2 N7 4.2876
R8 2 1 10g
.ends 
*******
.subckt 0603_744917130_30n 1 2
C1 1 N7 92.9835f
L1 1 N1 29.4n
L2 N1 N2 565.8118p
L3 N2 N3 1.0666n
L4 N3 N4 2.6552n
L5 N4 N5 81.2516p
L6 N5 N6 56.6032p
R1 2 N1 4.9144
R2 2 N2 1.5763
R3 2 N3 440.7233m
R4 2 N4 362.6318m
R5 2 N5 550.5651m
R6 2 N6 481.2351m
R7 2 N7 4.3357
R8 2 1 10g
.ends 
*******
.subckt 0603_744917133_33n 1 2
C1 1 N7 109.0794f
L1 1 N1 32.4n
L2 N1 N2 689.5176p
L3 N2 N3 1.3018n
L4 N3 N4 3.0957n
L5 N4 N5 83.3482p
L6 N5 N6 57.8621p
R1 2 N1 5.6981
R2 2 N2 1.7178
R3 2 N3 510.4188m
R4 2 N4 371.9058m
R5 2 N5 533.3970m
R6 2 N6 446.4882m
R7 2 N7 4.8651
R8 2 1 10g
.ends 
*******
.subckt 0603_744917136_36n 1 2
C1 1 N7 90.8914f
L1 1 N1 35.2n
L2 N1 N2 473.0414p
L3 N2 N3 1.3034n
L4 N3 N4 7.8780n
L5 N4 N5 136.7962p
L6 N5 N6 71.8756p
R1 2 N1 7.085
R2 2 N2 4.079
R3 2 N3 908.2290m
R4 2 N4 4.8542
R5 2 N5 1.2048
R6 2 N6 1.117
R7 2 N7 18.7415
R8 2 1 10g
.ends 
*******
.subckt 0603_744917139_39n 1 2
C1 1 N7 90.5148f
L1 1 N1 38.2n
L2 N1 N2 624.1302p
L3 N2 N3 1.0582n
L4 N3 N4 3.6988n
L5 N4 N5 97.2929p
L6 N5 N6 61.9433p
R1 2 N1 7.1253
R2 2 N2 4.1263
R3 2 N3 901.1808m
R4 2 N4 4.8037
R5 2 N5 347.5755m
R6 2 N6 892.6421m
R7 2 N7 11.7673
R8 2 1 10g
.ends 
*******
.subckt 0603_744917143_43n 1 2
C1 1 N7 90.8914f
L1 1 N1 41.5n
L2 N1 N2 775.7416p
L3 N2 N3 1.2813n
L4 N3 N4 6.0855n
L5 N4 N5 117.2872p
L6 N5 N6 66.9283p
R1 2 N1 6.0344
R2 2 N2 3.7764
R3 2 N3 901.1808m
R4 2 N4 4.8043
R5 2 N5 821.1040m
R6 2 N6 503.9431m
R7 2 N7 12.605
R8 2 1 10g
.ends 
*******
.subckt 0603_744917147_47n 1 2
C1 1 N7 80.9857f
L1 1 N1 45.5n
L2 N1 N2 968.6038p
L3 N2 N3 1.6047n
L4 N3 N4 11.6605n
L5 N4 N5 159.0036p
L6 N5 N6 66.8998p
R1 2 N1 7.0323
R2 2 N2 3.5204
R3 2 N3 3.4532
R4 2 N4 4.8129
R5 2 N5 1.0579
R6 2 N6 934.4013m
R7 2 N7 15.4871
R8 2 1 10g
.ends 
*******
.subckt 0603_744917151_51n 1 2
C1 1 N7 77.1684f
L1 1 N1 48n
L2 N1 N2 1.0920n
L3 N2 N3 690.7057p
L4 N3 N4 2.6906n
L5 N4 N5 104.1348p
L6 N5 N6 66.6695p
R1 2 N1 5.9609
R2 2 N2 3.1951
R3 2 N3 3.0625
R4 2 N4 4.813
R5 2 N5 1.079
R6 2 N6 968.0781m
R7 2 N7 15.7226
R8 2 1 10g
.ends 
*******
.subckt 0603_744917156_56n 1 2
C1 1 N7 73.3917f
L1 1 N1 53.5n
L2 N1 N2 1.3369n
L3 N2 N3 550.3818p
L4 N3 N4 3.3775n
L5 N4 N5 181.4284p
L6 N5 N6 67.1928p
R1 2 N1 5.7364
R2 2 N2 2.7623
R3 2 N3 2.5094
R4 2 N4 4.7957
R5 2 N5 636.8563m
R6 2 N6 296.1908m
R7 2 N7 16.6597
R8 2 1 10g
.ends 
*******
.subckt 0603_744917168_68n 1 2
C1 1 N7 70.4521f
L1 1 N1 65.5n
L2 N1 N2 2.2634n
L3 N2 N3 1.8432n
L4 N3 N4 7.1619n
L5 N4 N5 207.0687p
L6 N5 N6 67.0281p
R1 2 N1 6.0088
R2 2 N2 2.6481
R3 2 N3 2.4856
R4 2 N4 4.8018
R5 2 N5 898.3166m
R6 2 N6 814.6576m
R7 2 N7 19.4106
R8 2 1 10g
.ends 
*******
.subckt 0603_744917172_72n 1 2
C1 1 N7 75.0031f
L1 1 N1 69.5n
L2 N1 N2 2.5470n
L3 N2 N3 201.5151p
L4 N3 N4 5.2962n
L5 N4 N5 170.5809p
L6 N5 N6 66.3594p
R1 2 N1 6.3293
R2 2 N2 2.635
R3 2 N3 2.4566
R4 2 N4 4.7971
R5 2 N5 778.1208m
R6 2 N6 665.7349m
R7 2 N7 23.586
R8 2 1 10g
.ends 
*******
.subckt 0603_744917175_75n 1 2
C1 1 N7 75.0031f
L1 1 N1 72.5n
L2 N1 N2 2.5470n
L3 N2 N3 201.5151p
L4 N3 N4 5.2962n
L5 N4 N5 170.5809p
L6 N5 N6 66.3594p
R1 2 N1 6.3293
R2 2 N2 2.635
R3 2 N3 2.4566
R4 2 N4 4.7971
R5 2 N5 778.1208m
R6 2 N6 665.7349m
R7 2 N7 23.586
R8 2 1 10g
.ends 
*******
.subckt 0603_744917182_82n 1 2
C1 1 N7 70.4080f
L1 1 N1 79.5n
L2 N1 N2 2.9707n
L3 N2 N3 949.0093p
L4 N3 N4 5.5394n
L5 N4 N5 162.4296p
L6 N5 N6 66.0661p
R1 2 N1 6.6587
R2 2 N2 2.6694
R3 2 N3 2.4575
R4 2 N4 4.7981
R5 2 N5 824.0405m
R6 2 N6 727.0751m
R7 2 N7 26.5577
R8 2 1 10g
.ends 
*******
.subckt 0603_744917191_91n 1 2
C1 1 N7 65.0031f
L1 1 N1 88.5n
L2 N1 N2 2.9864n
L3 N2 N3 922.6129p
L4 N3 N4 4.7111n
L5 N4 N5 154.8249p
L6 N5 N6 66.0295p
R1 2 N1 6.6855
R2 2 N2 2.6751
R3 2 N3 2.4615
R4 2 N4 4.7976
R5 2 N5 808.8122m
R6 2 N6 707.7853m
R7 2 N7 26.921
R8 2 1 10g
.ends 
*******
.subckt 0603_744917210_100n 1 2
C1 1 N7 57.8827f
L1 1 N1 97n
L2 N1 N2 3.5296n
L3 N2 N3 6.4836n
L4 N3 N4 11.4964n
L5 N4 N5 210.3817p
L6 N5 N6 66.0670p
R1 2 N1 7.1589
R2 2 N2 2.3505
R3 2 N3 2.4747
R4 2 N4 4.8184
R5 2 N5 1.2793
R6 2 N6 1.249
R7 2 N7 30.4081
R8 2 1 10g
.ends 
*******
.subckt 0603_744917211_110n 1 2
C1 1 N7 60.9231f
L1 1 N1 107n
L2 N1 N2 4.1270n
L3 N2 N3 3.0107n
L4 N3 N4 5.8202n
L5 N4 N5 147.4963p
L6 N5 N6 65.4090p
R1 2 N1 7.6623
R2 2 N2 2.3617
R3 2 N3 2.3384
R4 2 N4 4.8111
R5 2 N5 1.1859
R6 2 N6 1.1521
R7 2 N7 33.9069
R8 2 1 10g
.ends 
*******
.subckt 0603_744917212_120n 1 2
C1 1 N7 60.0573f
L1 1 N1 117n
L2 N1 N2 4.6821n
L3 N2 N3 1.3148n
L4 N3 N4 11.6281n
L5 N4 N5 195.9287p
L6 N5 N6 65.5524p
R1 2 N1 8.4326
R2 2 N2 4.1154
R3 2 N3 4.43
R4 2 N4 4.851
R5 2 N5 2.6281
R6 2 N6 1.6584
R7 2 N7 36.4833
R8 2 1 10g
.ends 
*******
.subckt 0603_744917215_150n 1 2
C1 1 N7 57.8075f
L1 1 N1 146n
L2 N1 N2 5.6958n
L3 N2 N3 1.9155n
L4 N3 N4 10.5411n
L5 N4 N5 190.7349p
L6 N5 N6 65.5531p
R1 2 N1 9.3993
R2 2 N2 4.1626
R3 2 N3 4.4122
R4 2 N4 4.8629
R5 2 N5 2.6686
R6 2 N6 1.7561
R7 2 N7 40.8829
R8 2 1 10g
.ends 
*******
.subckt 0603_744917218_180n 1 2
C1 1 N7 54.9316f
L1 1 N1 175n
L2 N1 N2 6.3348n
L3 N2 N3 1.5278n
L4 N3 N4 19.8204n
L5 N4 N5 351.0641p
L6 N5 N6 69.4470p
R1 2 N1 13.2469
R2 2 N2 7.2671
R3 2 N3 6.5172
R4 2 N4 5.0279
R5 2 N5 4.1424
R6 2 N6 3.6105
R7 2 N7 55.7177
R8 2 1 10g
.ends 
*******
.subckt 0603_744917220_200n 1 2
C1 1 N7 48.4970f
L1 1 N1 194n
L2 N1 N2 7.3158n
L3 N2 N3 396.8938p
L4 N3 N4 16.9620n
L5 N4 N5 337.7420p
L6 N5 N6 69.4288p
R1 2 N1 13.7889
R2 2 N2 7.3409
R3 2 N3 6.4236
R4 2 N4 5.1023
R5 2 N5 4.252
R6 2 N6 3.7533
R7 2 N7 56.7415
R8 2 1 10g
.ends 
*******
.subckt 0603_744917221_210n 1 2
C1 1 N7 58.9094f
L1 1 N1 203n
L2 N1 N2 7.3572n
L3 N2 N3 1.7506n
L4 N3 N4 16.9596n
L5 N4 N5 337.7784p
L6 N5 N6 69.4315p
R1 2 N1 13.8002
R2 2 N2 7.3491
R3 2 N3 6.4306
R4 2 N4 5.1042
R5 2 N5 4.2547
R6 2 N6 3.7568
R7 2 N7 56.7817
R8 2 1 10g
.ends 
*******
.subckt 0603_744917222_220n 1 2
C1 1 N7 64.5788f
L1 1 N1 212n
L2 N1 N2 7.7293n
L3 N2 N3 5.1515n
L4 N3 N4 30.1566n
L5 N4 N5 418.3024p
L6 N5 N6 70.0959p
R1 2 N1 14.8058
R2 2 N2 7.5707
R3 2 N3 6.3644
R4 2 N4 5.4976
R5 2 N5 4.7995
R6 2 N6 4.4348
R7 2 N7 58.1716
R8 2 1 10g
.ends 
*******
.subckt 0603_744917225_250n 1 2
C1 1 N7 62.7154f
L1 1 N1 241n
L2 N1 N2 9.0536n
L3 N2 N3 14.9760n
L4 N3 N4 167.6496n
L5 N4 N5 427.4827p
L6 N5 N6 70.2568p
R1 2 N1 20.1725
R2 2 N2 7.8556
R3 2 N3 6.7206
R4 2 N4 5.5304
R5 2 N5 4.8419
R6 2 N6 4.4843
R7 2 N7 58.5371
R8 2 1 10g
.ends 
*******
.subckt 0603_744917227_270n 1 2
C1 1 N7 51.1909f
L1 1 N1 260n
L2 N1 N2 8.9284n
L3 N2 N3 9.7349n
L4 N3 N4 165.4156n
L5 N4 N5 426.6680p
L6 N5 N6 70.2126p
R1 2 N1 20.2728
R2 2 N2 7.5892
R3 2 N3 6.5038
R4 2 N4 5.5345
R5 2 N5 4.8472
R6 2 N6 4.4905
R7 2 N7 58.5809
R8 2 1 10g
.ends 
*******
.subckt 0603_744917230_300n 1 2
C1 1 N7 51.9731f
L1 1 N1 288n
L2 N1 N2 10.6836n
L3 N2 N3 9.9721n
L4 N3 N4 165.7836n
L5 N4 N5 426.3779p
L6 N5 N6 70.1938p
R1 2 N1 20.779
R2 2 N2 7.5846
R3 2 N3 6.4866
R4 2 N4 5.5353
R5 2 N5 4.8483
R6 2 N6 4.4918
R7 2 N7 58.6385
R8 2 1 10g
.ends 
*******
.subckt 0603_744917233_330n 1 2
C1 1 N7 51.3924f
L1 1 N1 317n
L2 N1 N2 10.7890n
L3 N2 N3 8.1173n
L4 N3 N4 170.9662n
L5 N4 N5 426.5206p
L6 N5 N6 70.1857p
R1 2 N1 22.2997
R2 2 N2 10.5158
R3 2 N3 9.4211
R4 2 N4 8.5392
R5 2 N5 6.854
R6 2 N6 5.5004
R7 2 N7 58.7808
R8 2 1 10g
.ends 
*******
.subckt 0603_744917236_360n 1 2
C1 1 N7 49.5965f
L1 1 N1 346n
L2 N1 N2 13.2037n
L3 N2 N3 8.7099n
L4 N3 N4 171.4330n
L5 N4 N5 426.9321p
L6 N5 N6 70.2092p
R1 2 N1 22.7224
R2 2 N2 10.5265
R3 2 N3 9.4227
R4 2 N4 8.5395
R5 2 N5 6.8546
R6 2 N6 5.5013
R7 2 N7 58.7865
R8 2 1 10g
.ends 
*******
.subckt 0603_744917239_390n 1 2
C1 1 N7 46.1100f
L1 1 N1 375n
L2 N1 N2 14.3011n
L3 N2 N3 10.8507n
L4 N3 N4 183.1007n
L5 N4 N5 427.9259p
L6 N5 N6 70.2332p
R1 2 N1 25.2993
R2 2 N2 14.5993
R3 2 N3 10.4974
R4 2 N4 10.543
R5 2 N5 8.8597
R6 2 N6 6.5097
R7 2 N7 68.8976
R8 2 1 10g
.ends 
*******
