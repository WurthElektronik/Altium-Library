**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT EMI Suppression Ferrite Bead (High Frequency) 
* Matchcode:              WE-CBF HF
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-30
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0402_742841160_600ohm 1 2
Rp 1 2 1567.537
Cp 1 2 0.101559359p
Rs 1 N3 0.82
L1 N3 2 0.660682809u
.ends 0402_742841160_600ohm
*******
.subckt 0402_742841210_1000ohm 1 2
Rp 1 2 1645.505
Cp 1 2 8.16284970000001E-02p
Rs 1 N3 0.9
L1 N3 2 1.422223u
.ends 0402_742841210_1000ohm
*******
.subckt 0402_742843122_220ohm 1 2
Rp 1 2 404.788433
Cp 1 2 0.154244614p
Rs 1 N3 0.25
L1 N3 2 0.341027576u
.ends 0402_742843122_220ohm
*******
.subckt 0603_742861118_180ohm 1 2
Rp 1 2 229.776461
Cp 1 2 0.31745586p
Rs 1 N3 0.25
L1 N3 2 0.375409809u
.ends 0603_742861118_180ohm
*******
.subckt 0603_742861160_600ohm 1 2
Rp 1 2 749.834927
Cp 1 2 0.159600804999999p
Rs 1 N3 0.27
L1 N3 2 1.460486u
.ends 0603_742861160_600ohm
*******
.subckt 0603_742861210_1000ohm 1 2
Rp 1 2 2431.131
Cp 1 2 0.093086003p
Rs 1 N3 1.2
L1 N3 2 1.270128u
.ends 0603_742861210_1000ohm
*******
.subckt 0603_742862160_600ohm 1 2
Rp 1 2 1431.286
Cp 1 2 0.121191332p
Rs 1 N3 0.8
L1 N3 2 0.719111746u
.ends 0603_742862160_600ohm
*******
.subckt 0603_742863122_220ohm 1 2
Rp 1 2 425.662883
Cp 1 2 0.184055236p
Rs 1 N3 0.13
L1 N3 2 0.35233079u
.ends 0603_742863122_220ohm
*******
.subckt 0603_742863147_470ohm 1 2
Rp 1 2 1038.428
Cp 1 2 0.095275095p
Rs 1 N3 0.19
L1 N3 2 0.823876562u
.ends 0603_742863147_470ohm
*******
.subckt 0603_742863160_600ohm 1 2
Rp 1 2 977.275205
Cp 1 2 0.139110959p
Rs 1 N3 0.22
L1 N3 2 0.620177887u
.ends 0603_742863160_600ohm
*******
