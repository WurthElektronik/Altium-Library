**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Film Capacitors
* Matchcode:             WCAP-FTX2
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 890324022007_15nF 1 2
Rser 1 3 0.129
Lser 2 4 0.000000003657
C1 3 4 0.000000015
Rpar 3 4 30000000000
.ends 890324022007_15nF
*******
.subckt 890324022007CS_15nF 1 2
Rser 1 3 0.129
Lser 2 4 0.000000003657
C1 3 4 0.000000015
Rpar 3 4 30000000000
.ends 890324022007CS_15nF
*******
.subckt 890324022017_68nF 1 2
Rser 1 3 0.081
Lser 2 4 0.000000005101
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890324022017_68nF
*******
.subckt 890324022017CS_68nF 1 2
Rser 1 3 0.081
Lser 2 4 0.000000005101
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890324022017CS_68nF
*******
.subckt 890324023002_5.6nF 1 2
Rser 1 3 0.181
Lser 2 4 0.000000007973
C1 3 4 0.0000000056
Rpar 3 4 30000000000
.ends 890324023002_5.6nF
*******
.subckt 890324023002CS_5.6nF 1 2
Rser 1 3 0.181
Lser 2 4 0.000000007973
C1 3 4 0.0000000056
Rpar 3 4 30000000000
.ends 890324023002CS_5.6nF
*******
.subckt 890324023003_6.8nF 1 2
Rser 1 3 0.165
Lser 2 4 0.000000005817
C1 3 4 0.0000000068
Rpar 3 4 30000000000
.ends 890324023003_6.8nF
*******
.subckt 890324023003CS_6.8nF 1 2
Rser 1 3 0.165
Lser 2 4 0.000000005817
C1 3 4 0.0000000068
Rpar 3 4 30000000000
.ends 890324023003CS_6.8nF
*******
.subckt 890324023004_8.2nF 1 2
Rser 1 3 0.136
Lser 2 4 0.000000006165
C1 3 4 0.0000000082
Rpar 3 4 30000000000
.ends 890324023004_8.2nF
*******
.subckt 890324023004CS_8.2nF 1 2
Rser 1 3 0.136
Lser 2 4 0.000000006165
C1 3 4 0.0000000082
Rpar 3 4 30000000000
.ends 890324023004CS_8.2nF
*******
.subckt 890324023006_10nF 1 2
Rser 1 3 0.135
Lser 2 4 0.000000006652
C1 3 4 0.00000001
Rpar 3 4 30000000000
.ends 890324023006_10nF
*******
.subckt 890324023006CS_10nF 1 2
Rser 1 3 0.135
Lser 2 4 0.000000006652
C1 3 4 0.00000001
Rpar 3 4 30000000000
.ends 890324023006CS_10nF
*******
.subckt 890324023007_12nF 1 2
Rser 1 3 0.152
Lser 2 4 0.000000007508
C1 3 4 0.000000012
Rpar 3 4 30000000000
.ends 890324023007_12nF
*******
.subckt 890324023007CS_12nF 1 2
Rser 1 3 0.152
Lser 2 4 0.000000007508
C1 3 4 0.000000012
Rpar 3 4 30000000000
.ends 890324023007CS_12nF
*******
.subckt 890324023008_15nF 1 2
Rser 1 3 0.13
Lser 2 4 0.00000000435
C1 3 4 0.000000015
Rpar 3 4 30000000000
.ends 890324023008_15nF
*******
.subckt 890324023008CS_15nF 1 2
Rser 1 3 0.13
Lser 2 4 0.00000000435
C1 3 4 0.000000015
Rpar 3 4 30000000000
.ends 890324023008CS_15nF
*******
.subckt 890324023010_18nF 1 2
Rser 1 3 0.0858385945068
Lser 2 4 8.0360172E-09
C1 3 4 0.000000018
Rpar 3 4 30000000000
.ends 890324023010_18nF
*******
.subckt 890324023010CS_18nF 1 2
Rser 1 3 0.198
Lser 2 4 0.000000012
C1 3 4 0.000000018
Rpar 3 4 30000000000
.ends 890324023010CS_18nF
*******
.subckt 890324023011_22nF 1 2
Rser 1 3 0.115
Lser 2 4 0.000000004093
C1 3 4 0.000000022
Rpar 3 4 30000000000
.ends 890324023011_22nF
*******
.subckt 890324023011CS_22nF 1 2
Rser 1 3 0.115
Lser 2 4 0.000000004093
C1 3 4 0.000000022
Rpar 3 4 30000000000
.ends 890324023011CS_22nF
*******
.subckt 890324023015_47nF 1 2
Rser 1 3 0.065
Lser 2 4 7.800475252E-09
C1 3 4 0.000000047
Rpar 3 4 30000000000
.ends 890324023015_47nF
*******
.subckt 890324023015CS_47nF 1 2
Rser 1 3 0.084
Lser 2 4 0.000000004714
C1 3 4 0.000000047
Rpar 3 4 30000000000
.ends 890324023015CS_47nF
*******
.subckt 890324023017_56nF 1 2
Rser 1 3 0.093
Lser 2 4 0.000000003499
C1 3 4 0.000000056
Rpar 3 4 30000000000
.ends 890324023017_56nF
*******
.subckt 890324023017CS_56nF 1 2
Rser 1 3 0.093
Lser 2 4 0.000000003499
C1 3 4 0.000000056
Rpar 3 4 30000000000
.ends 890324023017CS_56nF
*******
.subckt 890324023019_68nF 1 2
Rser 1 3 0.129
Lser 2 4 0.000000004657
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890324023019_68nF
*******
.subckt 890324023019CS_68nF 1 2
Rser 1 3 0.129
Lser 2 4 0.000000004657
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890324023019CS_68nF
*******
.subckt 890324023021_82nF 1 2
Rser 1 3 0.08
Lser 2 4 0.000000004262
C1 3 4 0.000000082
Rpar 3 4 30000000000
.ends 890324023021_82nF
*******
.subckt 890324023021CS_82nF 1 2
Rser 1 3 0.08
Lser 2 4 0.000000004262
C1 3 4 0.000000082
Rpar 3 4 30000000000
.ends 890324023021CS_82nF
*******
.subckt 890324023023_100nF 1 2
Rser 1 3 0.068
Lser 2 4 0.000000005686
C1 3 4 0.0000001
Rpar 3 4 30000000000
.ends 890324023023_100nF
*******
.subckt 890324023023CS_100nF 1 2
Rser 1 3 0.068
Lser 2 4 0.000000005686
C1 3 4 0.0000001
Rpar 3 4 30000000000
.ends 890324023023CS_100nF
*******
.subckt 890324023024_120nF 1 2
Rser 1 3 0.076
Lser 2 4 0.000000003321
C1 3 4 0.00000012
Rpar 3 4 30000000000
.ends 890324023024_120nF
*******
.subckt 890324023024CS_120nF 1 2
Rser 1 3 0.076
Lser 2 4 0.000000003321
C1 3 4 0.00000012
Rpar 3 4 30000000000
.ends 890324023024CS_120nF
*******
.subckt 890324023025_150nF 1 2
Rser 1 3 0.06
Lser 2 4 0.000000004594
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890324023025_150nF
*******
.subckt 890324023025CS_150nF 1 2
Rser 1 3 0.06
Lser 2 4 0.000000004594
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890324023025CS_150nF
*******
.subckt 890324023028_220nF 1 2
Rser 1 3 0.058
Lser 2 4 0.000000008265
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890324023028_220nF
*******
.subckt 890324023028CS_220nF 1 2
Rser 1 3 0.058
Lser 2 4 0.000000008265
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890324023028CS_220nF
*******
.subckt 890324024001_150nF 1 2
Rser 1 3 0.071
Lser 2 4 0.000000008975
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890324024001_150nF
*******
.subckt 890324024001CS_150nF 1 2
Rser 1 3 0.071
Lser 2 4 0.000000008975
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890324024001CS_150nF
*******
.subckt 890324024002_220nF 1 2
Rser 1 3 0.055
Lser 2 4 0.000000004818
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890324024002_220nF
*******
.subckt 890324024002CS_220nF 1 2
Rser 1 3 0.055
Lser 2 4 0.000000004818
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890324024002CS_220nF
*******
.subckt 890324024003_330nF 1 2
Rser 1 3 0.051
Lser 2 4 0.000000004813
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890324024003_330nF
*******
.subckt 890324024003CS_330nF 1 2
Rser 1 3 0.051
Lser 2 4 0.000000004813
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890324024003CS_330nF
*******
.subckt 890324024005_470nF 1 2
Rser 1 3 0.041
Lser 2 4 0.000000008759
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890324024005_470nF
*******
.subckt 890324024005CS_470nF 1 2
Rser 1 3 0.041
Lser 2 4 0.000000008759
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890324024005CS_470nF
*******
.subckt 890324025004_27nF 1 2
Rser 1 3 0.124
Lser 2 4 0.000000005256
C1 3 4 0.000000027
Rpar 3 4 30000000000
.ends 890324025004_27nF
*******
.subckt 890324025004CS_27nF 1 2
Rser 1 3 0.124
Lser 2 4 0.000000005256
C1 3 4 0.000000027
Rpar 3 4 30000000000
.ends 890324025004CS_27nF
*******
.subckt 890324025006_33nF 1 2
Rser 1 3 0.129
Lser 2 4 0.000000006876
C1 3 4 0.000000033
Rpar 3 4 30000000000
.ends 890324025006_33nF
*******
.subckt 890324025006CS_33nF 1 2
Rser 1 3 0.129
Lser 2 4 0.000000006876
C1 3 4 0.000000033
Rpar 3 4 30000000000
.ends 890324025006CS_33nF
*******
.subckt 890324025007_39nF 1 2
Rser 1 3 0.114
Lser 2 4 0.000000005321
C1 3 4 0.000000039
Rpar 3 4 30000000000
.ends 890324025007_39nF
*******
.subckt 890324025007CS_39nF 1 2
Rser 1 3 0.114
Lser 2 4 0.000000005321
C1 3 4 0.000000039
Rpar 3 4 30000000000
.ends 890324025007CS_39nF
*******
.subckt 890324025009_47nF 1 2
Rser 1 3 0.115
Lser 2 4 0.000000007853
C1 3 4 0.000000047
Rpar 3 4 30000000000
.ends 890324025009_47nF
*******
.subckt 890324025009CS_47nF 1 2
Rser 1 3 0.115
Lser 2 4 0.000000007853
C1 3 4 0.000000047
Rpar 3 4 30000000000
.ends 890324025009CS_47nF
*******
.subckt 890324025011_56nF 1 2
Rser 1 3 0.096
Lser 2 4 0.000000005899
C1 3 4 0.000000056
Rpar 3 4 30000000000
.ends 890324025011_56nF
*******
.subckt 890324025011CS_56nF 1 2
Rser 1 3 0.096
Lser 2 4 0.000000005899
C1 3 4 0.000000056
Rpar 3 4 30000000000
.ends 890324025011CS_56nF
*******
.subckt 890324025013_68nF 1 2
Rser 1 3 0.079
Lser 2 4 0.000000005773
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890324025013_68nF
*******
.subckt 890324025013CS_68nF 1 2
Rser 1 3 0.079
Lser 2 4 0.000000005773
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890324025013CS_68nF
*******
.subckt 890324025015_82nF 1 2
Rser 1 3 0.076
Lser 2 4 0.000000005628
C1 3 4 0.000000082
Rpar 3 4 30000000000
.ends 890324025015_82nF
*******
.subckt 890324025015CS_82nF 1 2
Rser 1 3 0.076
Lser 2 4 0.000000005628
C1 3 4 0.000000082
Rpar 3 4 30000000000
.ends 890324025015CS_82nF
*******
.subckt 890324025017_100nF 1 2
Rser 1 3 0.072
Lser 2 4 0.000000004703
C1 3 4 0.0000001
Rpar 3 4 30000000000
.ends 890324025017_100nF
*******
.subckt 890324025017CS_100nF 1 2
Rser 1 3 0.072
Lser 2 4 0.000000004703
C1 3 4 0.0000001
Rpar 3 4 30000000000
.ends 890324025017CS_100nF
*******
.subckt 890324025020_120nF 1 2
Rser 1 3 0.043
Lser 2 4 0.000000006282
C1 3 4 0.00000012
Rpar 3 4 30000000000
.ends 890324025020_120nF
*******
.subckt 890324025020CS_120nF 1 2
Rser 1 3 0.043
Lser 2 4 0.000000006282
C1 3 4 0.00000012
Rpar 3 4 30000000000
.ends 890324025020CS_120nF
*******
.subckt 890324025022_150nF 1 2
Rser 1 3 0.064
Lser 2 4 0.000000005433
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890324025022_150nF
*******
.subckt 890324025022CS_150nF 1 2
Rser 1 3 0.064
Lser 2 4 0.000000005433
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890324025022CS_150nF
*******
.subckt 890324025025_180nF 1 2
Rser 1 3 0.061
Lser 2 4 0.000000006237
C1 3 4 0.00000018
Rpar 3 4 30000000000
.ends 890324025025_180nF
*******
.subckt 890324025025CS_180nF 1 2
Rser 1 3 0.061
Lser 2 4 0.000000006237
C1 3 4 0.00000018
Rpar 3 4 30000000000
.ends 890324025025CS_180nF
*******
.subckt 890324025027_220nF 1 2
Rser 1 3 0.057
Lser 2 4 0.000000005375
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890324025027_220nF
*******
.subckt 890324025027CS_220nF 1 2
Rser 1 3 0.057
Lser 2 4 0.000000005375
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890324025027CS_220nF
*******
.subckt 890324025031_270nF 1 2
Rser 1 3 0.038
Lser 2 4 0.000000005786
C1 3 4 0.00000027
Rpar 3 4 30000000000
.ends 890324025031_270nF
*******
.subckt 890324025031CS_270nF 1 2
Rser 1 3 0.038
Lser 2 4 0.000000005786
C1 3 4 0.00000027
Rpar 3 4 30000000000
.ends 890324025031CS_270nF
*******
.subckt 890324025034_330nF 1 2
Rser 1 3 0.066
Lser 2 4 0.000000006443
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890324025034_330nF
*******
.subckt 890324025034CS_330nF 1 2
Rser 1 3 0.066
Lser 2 4 0.000000006443
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890324025034CS_330nF
*******
.subckt 890324025039_470nF 1 2
Rser 1 3 0.037
Lser 2 4 0.000000005157
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890324025039_470nF
*******
.subckt 890324025039CS_470nF 1 2
Rser 1 3 0.037
Lser 2 4 0.000000005157
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890324025039CS_470nF
*******
.subckt 890324025043_560nF 1 2
Rser 1 3 0.078
Lser 2 4 0.000000007377
C1 3 4 0.00000056
Rpar 3 4 17857142857.1429
.ends 890324025043_560nF
*******
.subckt 890324025043CS_560nF 1 2
Rser 1 3 0.078
Lser 2 4 0.000000007377
C1 3 4 0.00000056
Rpar 3 4 17857142857.1429
.ends 890324025043CS_560nF
*******
.subckt 890324025045_680nF 1 2
Rser 1 3 0.04
Lser 2 4 9.692641615E-09
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890324025045_680nF
*******
.subckt 890324025045CS_680nF 1 2
Rser 1 3 0.03
Lser 2 4 0.000000003685
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890324025045CS_680nF
*******
.subckt 890324025047CS_820nF 1 2
Rser 1 3 0.06
Lser 2 4 0.000000014
C1 3 4 0.00000082
Rpar 3 4 12195121951.2195
.ends 890324025047CS_820nF
*******
.subckt 890324026003_220nF 1 2
Rser 1 3 0.069
Lser 2 4 0.000000010762
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890324026003_220nF
*******
.subckt 890324026003CS_220nF 1 2
Rser 1 3 0.069
Lser 2 4 0.000000010762
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890324026003CS_220nF
*******
.subckt 890324026007CS_330nF 1 2
Rser 1 3 0.0942681692678
Lser 2 4 1.0933931837E-08
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890324026007CS_330nF
*******
.subckt 890324026018_560nF 1 2
Rser 1 3 0.059
Lser 2 4 0.000000008177
C1 3 4 0.00000056
Rpar 3 4 17857142857.1429
.ends 890324026018_560nF
*******
.subckt 890324026018CS_560nF 1 2
Rser 1 3 0.059
Lser 2 4 0.000000008177
C1 3 4 0.00000056
Rpar 3 4 17857142857.1429
.ends 890324026018CS_560nF
*******
.subckt 890324026020_680nF 1 2
Rser 1 3 0.063
Lser 2 4 0.000000001199
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890324026020_680nF
*******
.subckt 890324026020CS_680nF 1 2
Rser 1 3 0.063
Lser 2 4 0.000000001199
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890324026020CS_680nF
*******
.subckt 890324026024_820nF 1 2
Rser 1 3 0.046
Lser 2 4 0.000000009104
C1 3 4 0.00000082
Rpar 3 4 12195121951.2195
.ends 890324026024_820nF
*******
.subckt 890324026024CS_820nF 1 2
Rser 1 3 0.046
Lser 2 4 0.000000009104
C1 3 4 0.00000082
Rpar 3 4 12195121951.2195
.ends 890324026024CS_820nF
*******
.subckt 890324026027_1uF 1 2
Rser 1 3 0.044
Lser 2 4 0.000000009842
C1 3 4 0.000001
Rpar 3 4 10000000000
.ends 890324026027_1uF
*******
.subckt 890324026027CS_1uF 1 2
Rser 1 3 0.044
Lser 2 4 0.000000009842
C1 3 4 0.000001
Rpar 3 4 10000000000
.ends 890324026027CS_1uF
*******
.subckt 890324026030_1.5uF 1 2
Rser 1 3 0.046
Lser 2 4 0.000000014416
C1 3 4 0.0000015
Rpar 3 4 6666666666.66667
.ends 890324026030_1.5uF
*******
.subckt 890324026030CS_1.5uF 1 2
Rser 1 3 0.046
Lser 2 4 0.000000014416
C1 3 4 0.0000015
Rpar 3 4 6666666666.66667
.ends 890324026030CS_1.5uF
*******
.subckt 890324026034_2.2uF 1 2
Rser 1 3 0.04
Lser 2 4 0.000000010658
C1 3 4 0.0000022
Rpar 3 4 4545454545.45455
.ends 890324026034_2.2uF
*******
.subckt 890324026034CS_2.2uF 1 2
Rser 1 3 0.04
Lser 2 4 0.000000010658
C1 3 4 0.0000022
Rpar 3 4 4545454545.45455
.ends 890324026034CS_2.2uF
*******
.subckt 890324027006_680nF 1 2
Rser 1 3 0.063
Lser 2 4 0.000000012215
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890324027006_680nF
*******
.subckt 890324027006CS_680nF 1 2
Rser 1 3 0.063
Lser 2 4 0.000000012215
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890324027006CS_680nF
*******
.subckt 890324027012_1.2uF 1 2
Rser 1 3 0.041
Lser 2 4 0.000000017256
C1 3 4 0.0000012
Rpar 3 4 8333333333.33333
.ends 890324027012_1.2uF
*******
.subckt 890324027012CS_1.2uF 1 2
Rser 1 3 0.041
Lser 2 4 0.000000017256
C1 3 4 0.0000012
Rpar 3 4 8333333333.33333
.ends 890324027012CS_1.2uF
*******
.subckt 890324027025_3.3uF 1 2
Rser 1 3 0.022
Lser 2 4 0.00000001046
C1 3 4 0.0000033
Rpar 3 4 3030303030.30303
.ends 890324027025_3.3uF
*******
.subckt 890324027025CS_3.3uF 1 2
Rser 1 3 0.022
Lser 2 4 0.00000001046
C1 3 4 0.0000033
Rpar 3 4 3030303030.30303
.ends 890324027025CS_3.3uF
*******
.subckt 890324027030CS_4.7uF 1 2
Rser 1 3 0.04
Lser 2 4 0.000000023
C1 3 4 0.0000047
Rpar 3 4 2127659574.46809
.ends 890324027030CS_4.7uF
*******
.subckt 890324028008_6.8uF 1 2
Rser 1 3 0.017
Lser 2 4 0.000000013001
C1 3 4 0.0000068
Rpar 3 4 1470588235.29412
.ends 890324028008_6.8uF
*******
.subckt 890324028008CS_6.8uF 1 2
Rser 1 3 0.017
Lser 2 4 0.000000013001
C1 3 4 0.0000068
Rpar 3 4 1470588235.29412
.ends 890324028008CS_6.8uF
*******
