**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Common Mode Power Line Choke 
* Matchcode:              WE-CMB HC 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-26
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt S_7448225007_0.7m  1  2  3  4
X1  1  2  3  4  CMBHC  PARAMS:
+  L1=385.38e-6
+  L2=60.35e-006
+  L3=92.47e-006
+  L4=80.22e-006
+  L5=18e-009
+  C1=2e-012
+  C2=1e-012
+  Rs1=2928
+  Rs2=837
+  Rs3=1193
+  Rs4=1278
+  Rs5=549
+  R2=0.11
+  dL3=200e-009
+  dC3=5.3e-012
+  dL4=4.01e-009
+  dC4=4.63e-012
+  dR3=0.48
+  dR4=2980
+  dR5=0.98
+  dR6=366
+  Rdc=15m
+  ck=4pF
.ends  S_7448225007_0.7m
*****
.subckt S_7448227005_0.45m  1  2  3  4
X1  1  2  3  4  CMBHC  PARAMS:
+  L1=208.89e-006
+  L2=40.29e-006
+  L3=50e-06
+  L4=50e-06
+  L5=125.26e-006
+  C1=9.80e-012
+  C2=1.87e-012
+  Rs1=1440
+  Rs2=1206
+  Rs3=254
+  Rs4=188
+  Rs5=1400
+  R2=0.054
+  dL3=140e-009
+  dC3=4.6e-012
+  dL4=4.11e-009
+  dC4=0.33e-012
+  dR3=0.48
+  dR4=2280
+  dR5=10
+  dR6=316
+  Rdc=10m
+  ck=4pF
.ends  S_7448227005_0.45m
***** 
.subckt S_7448229004_0.35m  1  2  3  4
X1  1  2  3  4  CMBHC  PARAMS:
+  L1=60u
+  L2=50u
+  L3=72u
+  L4=2.5u
+  L5=3.8n
+  C1=1.4p
+  C2=2.1p
+  Rs1=600
+  Rs2=500
+  Rs3=500
+  Rs4=.600
+  Rs5=200
+  R2=1.41
+  dL3=50n
+  dC3=3.5p
+  dL4=1.31n
+  dC4=1.03p
+  dR3=0.48
+  dR4=801
+  dR5=0.78
+  dR6=126
+  Rdc=7m
+  ck=4pF
.ends  S_7448229004_0.35m
*****
.subckt S_74482210002_0.175m  1  2  3  4
X1  1  2  3  4  CMBHC  PARAMS:
+  L1=38.89e-006
+  L2=20.29e-006
+  L3=1e-09
+  L4=1e-09
+  L5=105.26e-006
+  C1=2263.80e-015
+  C2=3.13e-012
+  Rs1=440
+  Rs2=206
+  Rs3=254
+  Rs4=188
+  Rs5=1200
+  R2=0.054
+  dL3=50e-009
+  dC3=3e-012
+  dL4=1.351e-009
+  dC4=1.43e-015
+  dR3=0.48
+  dR4=880
+  dR5=1.88
+  dR6=166
+  Rdc=4m
+  ck=4pF
.ends  S_74482210002_0.175m
 ******
.subckt S_7448228002_0.175m  1 2 3 4
X1  1  2  3  4  CMBHC1  PARAMS:
+ L3=130u
+ Rs3=700
+ C1=1.8p
+ R2=1
+ L5=77u
+ C2=44.1p
+ Rs5=830
+ Rs1=0.1k
+ Rs2=10
+ Rs4=1
+ Rdc=6m
+ L1=0.8p
+ L2=1p
+ L4=1p
+ dR5=100
+ ck=7.5p
+ dL4=2n
+ dL3=0.05u
+ dC3=10.1p
+ dC4=1.1p
+ dR3=2.5k
+ dR6=1.53k
+ dR4=0.2k
.ends
****
.subckt S_7448226404_0.35m  1 2 3 4
X1  1  2  3  4  CMBHC1  PARAMS:
+ L3=250u
+ Rs3=1800
+ C1=2.3p
+ R2=1
+ L5=130u
+ C2=32.1p
+ Rs5=1650
+ Rs1=0.1k
+ Rs2=10
+ Rs4=1
+ Rdc=10m
+ L1=0.8p
+ L2=1p
+ L4=1p
+ dR5=100
+ ck=8p
+ dL4=4.5n
+ dL3=0.09u
+ dC3=10.1p
+ dC4=0.1p
+ dR3=2.0k
+ dR6=1.0k
+ dR4=0.27k
.ends 
*****
.subckt CMBHC  1  2  3  4  PARAMS:
R_R9  N12325  3  {R2}
R_R8  N13265  N13287  {Rs4}
Kn_K6  L_L11  L_L12  
+  L_L13  L_L14  0.9999
R_R3  N12571  N12583  {Rs3}
R_R10  N13777  4  {R2}
C_C10  N13029  N12821  {ck}
R_R20  N13215  N13229  {dR4}
L_L11  N12821  N12295  {dL4}
R_R17  N12267  N12273  {dR3}
L_L8  N13265  N13287  {L4}
R_R7  N13287  N13305  {Rs3}
L_L9  N12295  N12307  {L5}
Kn_K4  L_L7  L_L8  1
R_R2  N12583  N12599  {Rs2}
Kn_K5  L_L9  L_L10  1
R_R16  N13229  N13249  {dR6}
Kn_K7  L_L15  L_L16
+  L_L17  L_L18  0.9999
C_C5  N12273  N12289  {dC4}
L_L6  N13287  N13305  {L3}
L_L7  N12307  N12571  {L4}
R_R6  N13305  N13319  {Rs2}
R_R21  1  N12257  {Rdc}
Kn_K3  L_L5  L_L6  1
L_L16  N12257  N12799  {dL3}
C_C8  N13215  N13741  {dC3}
L_L18  N13023  N13215  {dL3}
R_R1  N12599  3  {Rs1}
R_R13  N12289  N12295  {dR5}
L_L4  N13305  N13319  {L2}
L_L5  N12571  N12583  {L3}
R_R15  N13755  N13249  {dR5}
R_R5  N13319  4  {Rs1}
R_R18  N12257  N12273  {dR4}
Kn_K2  L_L3  L_L4  1
R_R19  N13741  N13229  {dR3}
L_L15  N12799  N12273  {dL3}
L_L17  N13229  N13023  {dL3}
L_L3  N12583  N12599  {L2}
R_R11  N12295  N12307  {Rs5}
L_L2  N13319  4  {L1}
C_C4  N13249  N13265  {C2}
L_L10  N13249  N13265  {L5}
Kn_K1  L_L1  L_L2  1
R_R14  N12273  N12295  {dR6}
C_C6  N13229  N13755  {dC4}
L_L12  N12273  N12821  {dL4}
L_L14  N13029  N13229  {dL4}
L_L1  N12599  3  {L1}
C_C1  N12307  N12325  {C1}
R_R12  N13249  N13265  {Rs5}
C_C2  N13265  N13777  {C1}
R_R22  2  N13215  {Rdc}
C_C9  N13023  N12799  {ck}
R_R4  N12307  N12571  {Rs4}
C_C3  N12295  N12307  {C2}
L_L13  N13249  N13029  {dL4}
C_C7  N12257  N12267  {dC3}  
.ends  CMBHC
*****
.subckt CMBHC1 1 2 3 4 PARAMS:
+ L3=130u
+ Rs3=700
+ C1=1.8p
+ R2=1
+ L5=77u
+ C2=44.1p
+ Rs5=830
+ Rs1=0.1k
+ Rs2=10
+ Rs4=1
+ Rdc=1m
+ L1=0.8p
+ L2=1p
+ L4=1p
+ dR5=100
+ ck=7.5p
+ dL4=2n
+ dL3=0.05u
+ dC3=10.1p
+ dC4=1.1p
+ dR3=2.5k
+ dR6=1.53k
+ dR4=0.2k
L5 N009 N008 {L3}
C3 N002 N001 {C1}
L1 4 N010 {L1}
L3 N010 N009 {L2}
L6 N015 N014 {L3}
C4 N024 N013 {C1}
L2 3 N016 {L1}
L4 N016 N015 {L2}
L8 N014 N013 {L4}
L7 N008 N001 {L4}
L9 N001 N007 {L5}
L10 N013 N021 {L5}
R1 N003 1 {Rdc}
R2 N005 N003 {dR4}
C1 N004 N003 {dC3}
L17 N011 N003 {dL3}
L18 N017 N018 {dL3}
C2 N011 N018 {ck}
R3 N005 N004 {dR3}
R4 N019 N022 {dR3}
C9 N022 N017 {dC3}
R5 N019 N017 {dR4}
L19 N005 N011 {dL3}
L20 N018 N019 {dL3}
R6 N017 2 {Rdc}
R8 N007 N005 {dR6}
C10 N006 N005 {dC4}
L13 N012 N005 {dL4}
L14 N019 N020 {dL4}
C11 N012 N020 {ck}
R9 N007 N006 {dR5}
R10 N021 N023 {dR5}
C12 N023 N019 {dC4}
R11 N021 N019 {dR6}
L15 N007 N012 {dL4}
L16 N020 N021 {dL4}
R7 N001 N007 {Rs5}
C5 N001 N007 {C2}
R12 N013 N021 {Rs5}
C6 N013 N021 {C2}
R13 N008 N001 {Rs4}
R14 N009 N008 {Rs3}
R15 N010 N009 {Rs2}
R16 4 N010 {Rs1}
R17 N014 N013 {Rs4}
R18 N015 N014 {Rs3}
R19 N016 N015 {Rs2}
R20 3 N016 {Rs1}
R21 4 N002 {R2}
R22 3 N024 {R2}
K3 L5 L6 1
K2 L3 L4 1
K1 L1 L2 1
K4 L7 L8 1
K5 L9  L10 1
K7 L17 L18 L19 L20 0.9999
K6 L13 L14 L15 L16 0.9999
.ends
****