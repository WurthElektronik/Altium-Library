**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  MLCCs - Multilayer Ceramic Chip Capacitors
* Matchcode:              WCAP-CSGP_6-3V
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/19/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0201_885012104004_10nF 1 2
Rser 1 3 0.0627
Lser 2 4 0.000000000218
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012104004_10nF
*******
.subckt 0201_885012104003_100nF 1 2
Rser 1 3 0.02829
Lser 2 4 0.00000000018
C1 3 4 0.0000001
Rpar 3 4 500000000
.ends 0201_885012104003_100nF
*******
.subckt 0201_885012104009_100nF 1 2
Rser 1 3 0.0337
Lser 2 4 0.00000000018
C1 3 4 0.0000001
Rpar 3 4 500000000
.ends 0201_885012104009_100nF
*******
.subckt 0201_885012104010_220nF 1 2
Rser 1 3 0.043
Lser 2 4 0.00000000021
C1 3 4 0.00000022
Rpar 3 4 200000000
.ends 0201_885012104010_220nF
*******
.subckt 0201_885012104011_1uF 1 2
Rser 1 3 0.0109
Lser 2 4 0.00000000023
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0201_885012104011_1uF
*******
.subckt 0402_885012105001_100nF 1 2
Rser 1 3 0.0306025790761
Lser 2 4 3.00070139E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0402_885012105001_100nF
*******
.subckt 0402_885012105002_220nF 1 2
Rser 1 3 0.0133971746954
Lser 2 4 3.17565902E-10
C1 3 4 0.00000022
Rpar 3 4 500000000
.ends 0402_885012105002_220nF
*******
.subckt 0402_885012105003_330nF 1 2
Rser 1 3 0.0127725917953
Lser 2 4 3.17985991E-10
C1 3 4 0.00000033
Rpar 3 4 300000000
.ends 0402_885012105003_330nF
*******
.subckt 0402_885012105004_470nF 1 2
Rser 1 3 0.0135620044546
Lser 2 4 2.89834924E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0402_885012105004_470nF
*******
.subckt 0402_885012105005_680nF 1 2
Rser 1 3 0.00866869355558
Lser 2 4 3.2312296E-10
C1 3 4 0.00000068
Rpar 3 4 200000000
.ends 0402_885012105005_680nF
*******
.subckt 0402_885012105006_1uF 1 2
Rser 1 3 0.0122136788791
Lser 2 4 3.38680925E-10
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0402_885012105006_1uF
*******
.subckt 0402_885012105007_2.2uF 1 2
Rser 1 3 0.00909909650012
Lser 2 4 3.49876612E-10
C1 3 4 0.0000022
Rpar 3 4 20000000
.ends 0402_885012105007_2.2uF
*******
.subckt 0402_885012105008_4.7uF 1 2
Rser 1 3 0.00453732146966
Lser 2 4 3.78498478E-10
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0402_885012105008_4.7uF
*******
.subckt 0402_885012105020_10uF 1 2
Rser 1 3 0.0058
Lser 2 4 0.0000000008
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0402_885012105020_10uF
*******
.subckt 0603_885012106001_470nF 1 2
Rser 1 3 0.00946787785536
Lser 2 4 2.50326617E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0603_885012106001_470nF
*******
.subckt 0603_885012106002_680nF 1 2
Rser 1 3 0.0104592893966
Lser 2 4 3.4734058E-10
C1 3 4 0.00000068
Rpar 3 4 200000000
.ends 0603_885012106002_680nF
*******
.subckt 0603_885012106003_1uF 1 2
Rser 1 3 0.00760558670624
Lser 2 4 3.54495768E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012106003_1uF
*******
.subckt 0603_885012106004_2.2uF 1 2
Rser 1 3 0.00652337052819
Lser 2 4 4.58001637E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0603_885012106004_2.2uF
*******
.subckt 0603_885012106005_4.7uF 1 2
Rser 1 3 0.00436564105168
Lser 2 4 5.20484374E-10
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0603_885012106005_4.7uF
*******
.subckt 0603_885012106006_10uF 1 2
Rser 1 3 0.00407641026021
Lser 2 4 4.16060333E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0603_885012106006_10uF
*******
.subckt 0603_885012206001_470nF 1 2
Rser 1 3 0.00945
Lser 2 4 0.00000000041822
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0603_885012206001_470nF
*******
.subckt 0603_885012206002_1uF 1 2
Rser 1 3 0.00781
Lser 2 4 0.00000000043943
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012206002_1uF
*******
.subckt 0603_885012106033_47uF 1 2
Rser 1 3 0.00455
Lser 2 4 0.0000000012598
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 0603_885012106033_47uF
*******
.subckt 0805_885012107001_2.2uF 1 2
Rser 1 3 0.00487002224398
Lser 2 4 2.50543345E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012107001_2.2uF
*******
.subckt 0805_885012107002_3.3uF 1 2
Rser 1 3 0.00453837206006
Lser 2 4 2.98091685E-10
C1 3 4 0.0000033
Rpar 3 4 30000000
.ends 0805_885012107002_3.3uF
*******
.subckt 0805_885012107003_4.7uF 1 2
Rser 1 3 0.00422571742874
Lser 2 4 2.56201535E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0805_885012107003_4.7uF
*******
.subckt 0805_885012107004_10uF 1 2
Rser 1 3 0.00320609856405
Lser 2 4 3.83098838E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 0805_885012107004_10uF
*******
.subckt 0805_885012107005_22uF 1 2
Rser 1 3 0.00282261758127
Lser 2 4 5.44199046E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 0805_885012107005_22uF
*******
.subckt 0805_885012107006_47uF 1 2
Rser 1 3 0.00246814753418
Lser 2 4 4.62831333E-10
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 0805_885012107006_47uF
*******
.subckt 0805_885012207001_2.2uF 1 2
Rser 1 3 0.00442275214815
Lser 2 4 2.37717125E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012207001_2.2uF
*******
.subckt 0805_885012207002_4.7uF 1 2
Rser 1 3 0.011
Lser 2 4 0.0000000007
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0805_885012207002_4.7uF
*******
.subckt 0805_885012207003_10uF 1 2
Rser 1 3 0.00336648172245
Lser 2 4 4.89291579E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0805_885012207003_10uF
*******
.subckt 1206_885012108001_4.7uF 1 2
Rser 1 3 0.00600320174513
Lser 2 4 5.14564007E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012108001_4.7uF
*******
.subckt 1206_885012108002_10uF 1 2
Rser 1 3 0.00340980665018
Lser 2 4 8.40328091E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012108002_10uF
*******
.subckt 1206_885012108003_22uF 1 2
Rser 1 3 0.003095358264
Lser 2 4 8.67209117E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1206_885012108003_22uF
*******
.subckt 1206_885012108004_47uF 1 2
Rser 1 3 0.00304958303174
Lser 2 4 8.27626832E-10
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1206_885012108004_47uF
*******
.subckt 1206_885012108005_100uF 1 2
Rser 1 3 0.00189819698397
Lser 2 4 0.0000000009
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 1206_885012108005_100uF
*******
.subckt 1206_885012208001_2.2uF 1 2
Rser 1 3 0.00708971442636
Lser 2 4 4.50708422E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 1206_885012208001_2.2uF
*******
.subckt 1206_885012208002_4.7uF 1 2
Rser 1 3 0.00380516684832
Lser 2 4 4.86025433E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012208002_4.7uF
*******
.subckt 1206_885012208003_10uF 1 2
Rser 1 3 0.00257769589302
Lser 2 4 7.50158848E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012208003_10uF
*******
.subckt 1210_885012109001_10uF 1 2
Rser 1 3 0.00236975905543
Lser 2 4 7.97405226E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1210_885012109001_10uF
*******
.subckt 1210_885012109002_22uF 1 2
Rser 1 3 0.00298875292394
Lser 2 4 0.0000000009
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1210_885012109002_22uF
*******
.subckt 1210_885012109003_47uF 1 2
Rser 1 3 0.0033888514929
Lser 2 4 1.535140948E-09
C1 3 4 0.000047
Rpar 3 4 2000000
.ends 1210_885012109003_47uF
*******
.subckt 1210_885012109004_100uF 1 2
Rser 1 3 0.00239801642091
Lser 2 4 0.0000000009
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 1210_885012109004_100uF
*******
