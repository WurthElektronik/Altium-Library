**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT High Current Inductor 
* Matchcode:              WE-LHMD 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1008_74434301008082_8.2u 1 2 3 4 
Rdc1 1 N1 32m
Rp1 1 4 4786
Cp1 1 4 24.714p
L1 N1 4 9.395u

Rdc2 2 N2 32m
Rp2 2 3 4786
Cp2 2 3 24.714p
L2 N2 3 9.395u

Rg1 1 0 100meg
Rg2 2 0 100meg
Rg3 3 0 100meg
Rg4 4 0 100meg
.ends 1008_74434301008082_8.2u
******
.subckt 1008_74434301008100_10u 1 2 3 4
Rdc1 1 N1 45m
Rp1 1 4 4842
Cp1 1 4 28.715p
L1 N1 4 10.382u

Rdc2 2 N2 45m
Rp2 2 3 4842
Cp2 2 3 28.715p
L2 N2 3 10.382u
Rg1 1 0 100meg
Rg2 2 0 100meg
Rg3 3 0 100meg
Rg4 4 0 100meg
.ends 1008_74434301008100_10u
******
.subckt 1008_74434301008150_15u 1 2 3 4
Rdc1 1 N1 65m
Rp1 1 4 6736
Cp1 1 4 31.878p
L1 N1 4 16.8u

Rdc2 2 N2 65m
Rp2 2 3 6736
Cp2 2 3 31.878p
L2 N2 3 16.8u
Rg1 1 0 100meg
Rg2 2 0 100meg
Rg3 3 0 100meg
Rg4 4 0 100meg
.ends 1008_74434301008150_15u
******
.subckt 1008_74434301008220_22u 1 2 3 4
Rdc1 1 N1 105m
Rp1 1 4 5961
Cp1 1 4 27.708p
L1 N1 4 24.587u

Rdc2 2 N2 105m
Rp2 2 3 5961
Cp2 2 3 27.708p
L2 N2 3 24.587u
Rg1 1 0 100meg
Rg2 2 0 100meg
Rg3 3 0 100meg
Rg4 4 0 100meg
.ends 1008_74434301008220_22u
******
.subckt 1213_74434301213082_8.2u 1 2 3 4
Rdc1 1 N1 16m
Rp1 1 4 2383
Cp1 1 4 36.728p
L1 N1 4 9.245u

Rdc2 2 N2 16m
Rp2 2 3 2383
Cp2 2 3 36.728p
L2 N2 3 9.245u
Rg1 1 0 100meg
Rg2 2 0 100meg
Rg3 3 0 100meg
Rg4 4 0 100meg
.ends 1213_74434301213082_8.2u
******
.subckt 1213_74434301213100_10u 1 2 3 4
Rdc1 1 N1 20.5m
Rp1 1 4 2117
Cp1 1 4 37.603p
L1 N1 4 10.762u

Rdc2 2 N2 20.5m
Rp2 2 3 2117
Cp2 2 3 37.603p
L2 N2 3 10.762u
Rg1 1 0 100meg
Rg2 2 0 100meg
Rg3 3 0 100meg
Rg4 4 0 100meg
.ends 1213_74434301213100_10u
******
.subckt 1213_74434301213150_15u 1 2 3 4
Rdc1 1 N1 33.2m
Rp1 1 4 2122
Cp1 1 4 43.189p
L1 N1 4 16.33u

Rdc2 2 N2 33.2m
Rp2 2 3 2122
Cp2 2 3 43.189p
L2 N2 3 16.33u
Rg1 1 0 100meg
Rg2 2 0 100meg
Rg3 3 0 100meg
Rg4 4 0 100meg
.ends 1213_74434301213150_15u
******
.subckt 1213_74434301213220_22u 1 2 3 4
Rdc1 1 N1 50m
Rp1 1 4 4301
Cp1 1 4 40.517p
L1 N1 4 23.319u

Rdc2 2 N2 50m
Rp2 2 3 4301
Cp2 2 3 40.517p
L2 N2 3 23.319u
Rg1 1 0 100meg
Rg2 2 0 100meg
Rg3 3 0 100meg
Rg4 4 0 100meg
.ends 1213_74434301213220_22u
******
