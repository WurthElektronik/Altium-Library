**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Coupled Flatwire Inductor
* Matchcode:              WE-CFWI
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-17
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1310_74485540080_0.8u  1  2  3  4  PARAMS:
+  Cww=108p
+  Rp1=705.4
+  Cp1=2.628p
+  Lp1=0.908u
+  Rp2=705.4
+  Cp2=2.628p
+  Lp2=0.908u
+  RDC1=0.0016
+  RDC2=0.0016
+  K=0.925337776166087
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1310_74485540120_1.2u  1  2  3  4  PARAMS:
+  Cww=223p
+  Rp1=960.7
+  Cp1=3.927p
+  Lp1=1.261u
+  Rp2=960.7
+  Cp2=3.927p
+  Lp2=1.261u
+  RDC1=0.0024
+  RDC2=0.0024
+  K=0.944722181384559
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1310_74485540170_1.7u  1  2  3  4  PARAMS:
+  Cww=254p
+  Rp1=1234
+  Cp1=3.572p
+  Lp1=1.659u
+  Rp2=1234
+  Cp2=3.572p
+  Lp2=1.659u
+  RDC1=0.0033
+  RDC2=0.0033
+  K=0.958859616787506
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1310_74485540220_2.2u  1  2  3  4  PARAMS:
+  Cww=279p
+  Rp1=1606
+  Cp1=3.806p
+  Lp1=2.279u
+  Rp2=1606
+  Cp2=3.806p
+  Lp2=2.279u
+  RDC1=0.0042
+  RDC2=0.0042
+  K=0.956793888700459
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1310_74485540290_2.9u  1  2  3  4  PARAMS:
+  Cww=384p
+  Rp1=2102
+  Cp1=3.772p
+  Lp1=2.772u
+  Rp2=2102
+  Cp2=3.772p
+  Lp2=2.772u
+  RDC1=0.0056
+  RDC2=0.0056
+  K=0.964543844304761
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1310_74485540350_3.5u  1  2  3  4  PARAMS:
+  Cww=417p
+  Rp1=2626
+  Cp1=3.533p
+  Lp1=3.53u
+  Rp2=2626
+  Cp2=3.533p
+  Lp2=3.53u
+  RDC1=0.0075
+  RDC2=0.0075
+  K=0.969241234899017
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1312_74485540680_6.8u  1  2  3  4  PARAMS:
+  Cww=556p
+  Rp1=4005
+  Cp1=4.764p
+  Lp1=6.508u
+  Rp2=4005
+  Cp2=4.764p
+  Lp2=6.508u
+  RDC1=0.0113
+  RDC2=0.0113
+  K=0.986154146165801
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1312_74485540820_8.2u  1  2  3  4  PARAMS:
+  Cww=573p
+  Rp1=5043
+  Cp1=4.715p
+  Lp1=9.462u
+  Rp2=5043
+  Cp2=4.715p
+  Lp2=9.462u
+  RDC1=0.013
+  RDC2=0.013
+  K=0.987420882906575
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1312_74485540101_10u  1  2  3  4  PARAMS:
+  Cww=684p
+  Rp1=5877
+  Cp1=4.596p
+  Lp1=9.706u
+  Rp2=5877
+  Cp2=4.596p
+  Lp2=9.706u
+  RDC1=0.0139
+  RDC2=0.0139
+  K=0.989141041510259
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1813_74485542680_6.8u  1  2  3  4  PARAMS:
+  Cww=549p
+  Rp1=3794
+  Cp1=6.578p
+  Lp1=6.782u
+  Rp2=3794
+  Cp2=6.578p
+  Lp2=6.782u
+  RDC1=0.0061
+  RDC2=0.0061
+  K=0.983541021603304
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1813_74485542820_8.2u  1  2  3  4  PARAMS:
+  Cww=645p
+  Rp1=6040
+  Cp1=7.414p
+  Lp1=8.521u
+  Rp2=6040
+  Cp2=7.414p
+  Lp2=8.521u
+  RDC1=0.0084
+  RDC2=0.0084
+  K=0.985875864149334
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1813_74485542101_10u  1  2  3  4  PARAMS:
+  Cww=767p
+  Rp1=7360
+  Cp1=6.196p
+  Lp1=10.196u
+  Rp2=7360
+  Cp2=6.196p
+  Lp2=10.196u
+  RDC1=0.011
+  RDC2=0.011
+  K=0.987420882906575
C_C1 3 1 {Cww/2}
R_R50 3 1 5000g
C_C2 2 4 {Cww/2}
C_C5 2 3 {Cp1}
R_R1 2 N05454 {RDC1}
R_R2 2 3 {Rp1}
L_L1 N05454 3 {Lp1}
L_L2 N05750 1 {Lp2}
C_C6 4 1 {Cp2}
R_R3 4 1 {Rp2}
R_R4 4 N05750 {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
