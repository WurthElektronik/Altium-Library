**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT Power Inductor
* Matchcode:             WE-LQFS
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/10/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 3818_74406032010_1u 1 2
Rp 1 2 1464.724593754
Cp 1 2 0.4433002p
Rs 1 N3 0.026
L1 N3 2 0.815049662u
.ends 3818_74406032010_1u
*******
.subckt 3818_74406032015_1.5u 1 2
Rp 1 2 1661.133174
Cp 1 2 0.488819396p
Rs 1 N3 0.032
L1 N3 2 1.209449053u
.ends 3818_74406032015_1.5u
*******
.subckt 3818_74406032033_3.3u 1 2
Rp 1 2 3688.21128
Cp 1 2 0.530944336p
Rs 1 N3 0.064
L1 N3 2 2.675333849u
.ends 3818_74406032033_3.3u
*******
.subckt 3818_74406032047_4.7u 1 2
Rp 1 2 5470.059477
Cp 1 2 0.572256871p
Rs 1 N3 0.092
L1 N3 2 4.445113865u
.ends 3818_74406032047_4.7u
*******
.subckt 3818_74406032068_6.8u 1 2
Rp 1 2 5237.842532
Cp 1 2 0.665779819p
Rs 1 N3 0.127
L1 N3 2 6.264793582u
.ends 3818_74406032068_6.8u
*******
.subckt 3818_74406032100_10u 1 2
Rp 1 2 6292.074873
Cp 1 2 0.714631779p
Rs 1 N3 0.19
L1 N3 2 9.293387986u
.ends 3818_74406032100_10u
*******
.subckt 3818_74406032220_22u 1 2
Rp 1 2 9156.93522
Cp 1 2 0.884349082p
Rs 1 N3 0.401
L1 N3 2 22.9186456u
.ends 3818_74406032220_22u
*******
.subckt 3818_74406032330_33u 1 2
Rp 1 2 10918.67563
Cp 1 2 0.852066811p
Rs 1 N3 0.596
L1 N3 2 33.96214681u
.ends 3818_74406032330_33u
*******
.subckt 3818_74406032470_47u 1 2
Rp 1 2 14593.16774
Cp 1 2 0.836838329p
Rs 1 N3 0.834
L1 N3 2 49.06231398u
.ends 3818_74406032470_47u
*******
.subckt 3818_74406032101_100u 1 2
Rp 1 2 50357.67723
Cp 1 2 0.812990187p
Rs 1 N3 2.064
L1 N3 2 105.9848158u
.ends 3818_74406032101_100u
*******
.subckt 4818_74406042010_1u 1 2
Rp 1 2 1274.36368248571
Cp 1 2 0.5312728290537p
Rs 1 N3 0.019
L1 N3 2 0.8543352847166u
.ends 4818_74406042010_1u
*******
.subckt 4818_74406042015_1.5u 1 2
Rp 1 2 1814.95268867905
Cp 1 2 0.624419061307p
Rs 1 N3 0.025
L1 N3 2 1.30135618449143u
.ends 4818_74406042015_1.5u
*******
.subckt 4818_74406042022_2.2u 1 2
Rp 1 2 2368.12860174742
Cp 1 2 0.7352803846252p
Rs 1 N3 0.033
L1 N3 2 1.95297608861u
.ends 4818_74406042022_2.2u
*******
.subckt 4818_74406042033_3.3u 1 2
Rp 1 2 4736.03585966
Cp 1 2 1.09931748233p
Rs 1 N3 0.051
L1 N3 2 2.6054895112u
.ends 4818_74406042033_3.3u
*******
.subckt 4818_74406042047_4.7u 1 2
Rp 1 2 4814.18474981356
Cp 1 2 0.746166238624889p
Rs 1 N3 0.058
L1 N3 2 4.28567924260445u
.ends 4818_74406042047_4.7u
*******
.subckt 4818_74406042068_6.8u 1 2
Rp 1 2 7621.84117173571
Cp 1 2 1.08546710655857p
Rs 1 N3 0.081
L1 N3 2 6.72210857973u
.ends 4818_74406042068_6.8u
*******
.subckt 4818_74406042100_10u 1 2
Rp 1 2 9185.87299047
Cp 1 2 1.269171230004p
Rs 1 N3 0.111
L1 N3 2 9.454964068034u
.ends 4818_74406042100_10u
*******
.subckt 4818_74406042220_22u 1 2
Rp 1 2 19600.30355055
Cp 1 2 1.2041750408p
Rs 1 N3 0.283
L1 N3 2 21.72285997065u
.ends 4818_74406042220_22u
*******
.subckt 4818_74406042330_33u 1 2
Rp 1 2 26452.5732648571
Cp 1 2 1.24415788557714p
Rs 1 N3 0.407
L1 N3 2 32.1265300643143u
.ends 4818_74406042330_33u
*******
.subckt 4818_74406042470_47u 1 2
Rp 1 2 36664.6087587625
Cp 1 2 1.26516702855125p
Rs 1 N3 0.523
L1 N3 2 47.6683177326875u
.ends 4818_74406042470_47u
*******
.subckt 4818_74406042101_100u 1 2
Rp 1 2 65622.8858187
Cp 1 2 1.06980957186167p
Rs 1 N3 1.155
L1 N3 2 101.7558628034u
.ends 4818_74406042101_100u
*******
.subckt 4828_74406043012_1.2u 1 2
Rp 1 2 1125.1398015622
Cp 1 2 0.474347597678p
Rs 1 N3 0.018
L1 N3 2 1.07198872518u
.ends 4828_74406043012_1.2u
*******
.subckt 4828_74406043027_2.7u 1 2
Rp 1 2 2488.14420625833
Cp 1 2 0.725892531447833p
Rs 1 N3 0.027
L1 N3 2 2.481477322245u
.ends 4828_74406043027_2.7u
*******
.subckt 4828_74406043047_4.7u 1 2
Rp 1 2 4281.01908565286
Cp 1 2 0.882774464673857p
Rs 1 N3 0.042
L1 N3 2 4.47098537522571u
.ends 4828_74406043047_4.7u
*******
.subckt 4828_74406043068_6.8u 1 2
Rp 1 2 5463.2556027975
Cp 1 2 1.00090833700263p
Rs 1 N3 0.053
L1 N3 2 6.11750429502375u
.ends 4828_74406043068_6.8u
*******
.subckt 4828_74406043100_10u 1 2
Rp 1 2 7707.73858963333
Cp 1 2 1.35466615639333p
Rs 1 N3 0.072
L1 N3 2 9.08862383167u
.ends 4828_74406043100_10u
*******
.subckt 4828_74406043220_22u 1 2
Rp 1 2 16379.99510914
Cp 1 2 1.701638601062p
Rs 1 N3 0.143
L1 N3 2 22.54494837468u
.ends 4828_74406043220_22u
*******
.subckt 4828_74406043330_33u 1 2
Rp 1 2 24424.54399654
Cp 1 2 1.766709646812p
Rs 1 N3 0.209
L1 N3 2 33.93591268674u
.ends 4828_74406043330_33u
*******
.subckt 4828_74406043470_47u 1 2
Rp 1 2 32033.7344681667
Cp 1 2 1.91601989032667p
Rs 1 N3 0.216
L1 N3 2 45.4291974366u
.ends 4828_74406043470_47u
*******
.subckt 4828_74406043101_100u 1 2
Rp 1 2 62354.5865286
Cp 1 2 2.20914984961667p
Rs 1 N3 0.5
L1 N3 2 92.2579742918667u
.ends 4828_74406043101_100u
*******
.subckt 4828_74406043221_220u 1 2
Rp 1 2 146886.232786889
Cp 1 2 2.01937777070222p
Rs 1 N3 1.105
L1 N3 2 238.836027727778u
.ends 4828_74406043221_220u
*******
.subckt 4828_74406043331_330u 1 2
Rp 1 2 204781.0899775
Cp 1 2 2.5023004055175p
Rs 1 N3 1.554
L1 N3 2 300.00291584625u
.ends 4828_74406043331_330u
*******
.subckt 4828_74406043471_470u 1 2
Rp 1 2 571274.328987125
Cp 1 2 2.51133918219375p
Rs 1 N3 2.336
L1 N3 2 441.429966329125u
.ends 4828_74406043471_470u
*******
