**************************************************
* Manufacturer:           Würth Elektronik 
* Kinds:                  Common Mode Line Filter 
* Matchcode:              WE-CNSA
* Library Type:           LTspice
* Version:                rev23a
* Created/modified by:    Ella      
* Date and Time:          2023-07-24
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2023 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0805_784231061_67ohm 1 2 3 4
X1  1  2  3  4  CNSA  
+  L1=61.3001n
+  L2=62.1620n
+  L3=13.3422n
+  L4=54.6785n
+  C1=35.2735p
+  RS1=97.7477
+  RS2=9.2767
+  RS3=824.2056
+  RS4=3.8468k
+  R2=715.7781
+  dL3=343.8576p
+  dC3=6.0134p
+  DR3=675.6842
+  DR4=142.9781
+  Rdc=0.25
+  ck=5.0910p
.ends 0805_784231061_67ohm
*****
.subckt 0805_784231091_90ohm 1 2 3 4
X1  1  2  3  4  CNSA  PARAMS:
+  L1=50.6597n
+  L2=95.1175n
+  L3=15.7910n
+  L4=6.7634n
+  C1=13.9595f
+  RS1=729.4963
+  RS2=156.2918
+  RS3=379.4377
+  RS4=410.0680
+  R2=325.2338
+  dL3=391.8602p
+  dC3=106.6866f
+  DR3=168.0690
+  DR4=359.5189
+  Rdc=0.3
+  ck=3.3772p
.ends 0805_784231091_90ohm
*****
.subckt 0805_784231121_120ohm 1 2 3 4
X1  1  2  3  4  CNSA  PARAMS:
+  L1=55.0197n
+  L2=70.4975n
+  L3=110.2943n
+  L4=48.3324n
+  C1=32.6036f
+  RS1=193.3394
+  RS2=28.5251
+  RS3=163.6962
+  RS4=783.7053
+  R2=35.2518
+  dL3=336.5622p
+  dC3=9.9999f
+  DR3=10.0005
+  DR4=149.1075
+  Rdc=0.3
+  ck=5.4036p
.ends 0805_784231121_120ohm
*****
.subckt 0805_784231181_180ohm 1 2 3 4
X1  1  2  3  4  CNSA  PARAMS:
+  L1=259.4568n
+  L2=52.8697n
+  L3=37.0959n
+  L4=42.4253n
+  C1=11.4100f
+  RS1=305.2461
+  RS2=389.6341
+  RS3=458.6012
+  RS4=543.3033
+  R2=20.0553
+  dL3=454.7764p
+  dC3=17.1002p
+  DR3=179.9805
+  DR4=518.5033
+  Rdc=0.35
+  ck=5.3204p
.ends 0805_784231181_180ohm
*****
.subckt 0805_784231261_260ohm 1 2 3 4
X1  1  2  3  4  CNSA  PARAMS:
+  L1=329.8253n
+  L2=74.0714n
+  L3=69.6330n
+  L4=68.6305n
+  C1=28.6298f
+  RS1=392.5062
+  RS2=626.6374
+  RS3=628.3177
+  RS4=620.2937
+  R2=12.8183
+  dL3=688.1120p
+  dC3=11.3829f
+  DR3=1.0002
+  DR4=287.7703
+  Rdc=0.4
+  ck=2.2307p
.ends 0805_784231261_260ohm
*****
.subckt 0805_784231371_370ohm 1 2 3 4
X1  1  2  3  4  CNSA  PARAMS:
+  L1=501.9526n
+  L2=107.6264n
+  L3=106.3904n
+  L4=106.1505n
+  C1=28.3149f
+  RS1=482.1618
+  RS2=730.1847
+  RS3=729.4588
+  RS4=729.6500
+  R2=13.7909
+  dL3=433.0409p
+  dC3=70.7123f
+  DR3=9.9765
+  DR4=123.3352
+  Rdc=0.45
+  ck=8.0772p
.ends 0805_784231371_370ohm
*****
.subckt 1210_784234101_100u 1 2 3 4
X1  1  2  3  4  CNSA1  PARAMS:
+ dL3=3.7524n
+ dL4=574.0956p
+ dC3=599.8144p
+ dC4=15.4698p
+ dR3=267.9220
+ dR4=90.0294
+ dR5=214.3516
+ dR6=229.9689
+ ck=17.6783p
+ L1=67.7625u
+ L2=97.4558n
+ L3=50.0240n
+ L4=20.0097n
+ L5=3.2345n
+ C1=79.6877f
+ C2=78.3484f
+ RS1=30.2592k
+ RS2=2.5000k
+ RS3=199.9976
+ RS4=199.9968
+ Rs5=1.4862
+ R2=99.9304
+ Rdc=3.36
.ends 1210_784234101_100u
*****
.subckt 1210_784234201_200u 1 2 3 4
X1  1  2  3  4  CNSA1  PARAMS:
+ dL3=6.0010n
+ dL4=717.6097p
+ dC3=599.5379p
+ dC4=15.1406p
+ dR3=267.8192
+ dR4=90.0148
+ dR5=104.3158
+ dR6=109.9709
+ ck=26.0743p
+ L1=144.3849u
+ L2=99.5775n
+ L3=50.0379n
+ L4=20.0425n
+ L5=3.2344n
+ C1=76.1033f
+ C2=78.3479f
+ RS1=60.5625k
+ RS2=2.5000k
+ RS3=200.0011
+ RS4=199.9991
+ Rs5=1.4862
+ R2=99.9304
+ Rdc=5.5
.ends 1210_784234201_200u
*****
.SUBCKT  CNSA1  1  2  3  4  PARAMS:
L5 N009 N008 {L3}
C3 N002 N001 {C1}
L1 3 N010 {L1}
L3 N010 N009 {L2}
L6 N015 N014 {L3}
C4 N024 N013 {C1}
L2 4 N016 {L1}
L4 N016 N015 {L2}
L8 N014 N013 {L4}
L7 N008 N001 {L4}
L9 N001 N007 {L5}
L10 N013 N021 {L5}
R1 N003 1 {Rdc}
R2 N005 N003 {dR4}
C1 N004 N003 {dC3}
L17 N011 N003 {dL3}
L18 N017 N018 {dL3}
C2 N011 N018 {ck}
R3 N005 N004 {dR3}
R4 N019 N022 {dR3}
C9 N022 N017 {dC3}
R5 N019 N017 {dR4}
L19 N005 N011 {dL3}
L20 N018 N019 {dL3}
R6 N017 2 {Rdc}
R8 N007 N005 {dR6}
C10 N006 N005 {dC4}
L13 N012 N005 {dL4}
L14 N019 N020 {dL4}
C11 N012 N020 {ck}
R9 N007 N006 {dR5}
R10 N021 N023 {dR5}
C12 N023 N019 {dC4}
R11 N021 N019 {dR6}
L15 N007 N012 {dL4}
L16 N020 N021 {dL4}
R7 N001 N007 {Rs5}
C5 N001 N007 {C2}
R12 N013 N021 {Rs5}
C6 N013 N021 {C2}
R13 N008 N001 {Rs4}
R14 N009 N008 {Rs3}
R15 N010 N009 {Rs2}
R16 3 N010 {Rs1}
R17 N014 N013 {Rs4}
R18 N015 N014 {Rs3}
R19 N016 N015 {Rs2}
R20 4 N016 {Rs1}
R21 3 N002 {R2}
R22 4 N024 {R2}
K3 L5 L6 1
K2 L3 L4 1
K1 L1 L2 1
K4 L7 L8 1
K5 L9  L10 1
K6_1 L13 L14 0.9999
K6_2 L13 L15 0.9999
K6_3 L13 L16 0.9999
K6_4 L14 L15 0.9999
K6_5 L14 L16 0.9999
K6_6 L15 L16 0.9999
K7_1 L17 L18 0.9999
K7_2 L17 L19 0.9999
K7_3 L17 L20 0.9999
K7_4 L18 L19 0.9999
K7_5 L18 L20 0.9999
K7_6 L19 L20 0.9999
.ends  CNSA1
*****
.SUBCKT  CNSA  1  2  3  4  PARAMS:
R_R47  N21893  N21911  {Rs3}
R_R43  N21425  N21441  {Rs2}
R_R4  N22217  N21871  {dR3}
L_L3  N21425  N21441  {L2}
L_L8  N21871  N21893  {L4}
Kn_K1  L_L1  L_L2  1
R_R37  N21241  3  {R2}
R_R48  N21911  N21925  {Rs2}
R_R44  N21441  3  {Rs1}
C_C4  N21871  N22231  {C1}
L_L1  N21441  3  {L1}
C_C1  N21207  N21217  {dC3}
L_L6  N21893  N21911  {L3}
R_R1  1  N21207  {Rdc}
L_L17  N21207  N21585  {dL3}
R_R49  N21925  4  {Rs1}
Kn_K5_1  L_L17  L_L18  0.9999
Kn_K5_2  L_L17  L_L19  0.9999
Kn_K5_3  L_L17  L_L20  0.9999
Kn_K5_4  L_L18  L_L19  0.9999
Kn_K5_5  L_L18  L_L20  0.9999
Kn_K5_6  L_L19  L_L20  0.9999
R_R3  N21217  N21223  {dR3}
R_R55  N22231  4  {R2}
L_L4  N21911  N21925  {L2}
R_R2  N21207  N21223  {dR4}
L_L19  N21585  N21223  {dL3}
R_R6  2  N21857  {Rdc}
C_C2  N21731  N21585  {ck}
Kn_K4  L_L7  L_L8  1
L_L2  N21925  4  {L1}
R_R41  N21223  N21413  {Rs4}
L_L7  N21223  N21413  {L4}
R_R5  N21857  N21871  {dR4}
L_L18  N21731  N21857  {dL3}
Kn_K3  L_L5  L_L6  1
R_R46  N21871  N21893  {Rs4}
R_R42  N21413  N21425  {Rs3}
L_L5  N21413  N21425  {L3}
C_C9  N21857  N22217  {dC3}
L_L20  N21871  N21731  {dL3}
Kn_K2  L_L3  L_L4  1
C_C3  N21223  N21241  {C1}
.ends  CNSA
*****