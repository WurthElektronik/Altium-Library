**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Multi-Turn Ratio coupled Inductor 
* Matchcode:              WE-MTCI 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 5030_744889015100_10u  1  2  3  4  PARAMS:
+  Cww=9.5p
+  Rp1=9168
+  Cp1=9.155p
+  Lp1=10u
+  Rp2=20761
+  Cp2=5.514p
+  Lp2=22.5u
+  RDC1=0.349
+  RDC2=0.408
+  K=0.992191737742481
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_744889020100_10u  1  2  3  4  PARAMS:
+  Cww=10.2p
+  Rp1=6032
+  Cp1=13.907p
+  Lp1=10u
+  Rp2=31099
+  Cp2=3.902p
+  Lp2=40u
+  RDC1=0.358
+  RDC2=0.552
+  K=0.993856126408647
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_744889030100_10u  1  2  3  4  PARAMS:
+  Cww=13.6p
+  Rp1=5042
+  Cp1=29.032p
+  Lp1=10u
+  Rp2=57172
+  Cp2=4.282p
+  Lp2=90u
+  RDC1=0.363
+  RDC2=0.846
+  K=0.996828303504002
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_744889015220_22u  1  2  3  4  PARAMS:
+  Cww=12.1p
+  Rp1=19692
+  Cp1=8.558p
+  Lp1=22u
+  Rp2=19477
+  Cp2=8.547p
+  Lp2=49.5u
+  RDC1=0.662
+  RDC2=0.874
+  K=0.993615985817825
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_744889020220_22u  1  2  3  4  PARAMS:
+  Cww=13.2p
+  Rp1=16198
+  Cp1=17.947p
+  Lp1=22u
+  Rp2=34255
+  Cp2=5.509p
+  Lp2=88u
+  RDC1=0.712
+  RDC2=1.208
+  K=0.99572951785476
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_744889030220_22u  1  2  3  4  PARAMS:
+  Cww=14.9p
+  Rp1=11548
+  Cp1=29.125p
+  Lp1=22u
+  Rp2=127841
+  Cp2=4.581p
+  Lp2=198u
+  RDC1=0.732
+  RDC2=1.872
+  K=0.997851226740274
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_744889015330_33u  1  2  3  4  PARAMS:
+  Cww=17.9p
+  Rp1=14271
+  Cp1=8.324p
+  Lp1=33u
+  Rp2=63698
+  Cp2=5.312p
+  Lp2=74.25u
+  RDC1=1.338
+  RDC2=1.782
+  K=0.995342690085717
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_744889020330_33u  1  2  3  4  PARAMS:
+  Cww=18.9p
+  Rp1=16972
+  Cp1=15.439p
+  Lp1=33u
+  Rp2=55012
+  Cp2=4.466p
+  Lp2=132u
+  RDC1=1.383
+  RDC2=2.418
+  K=0.996775103050134
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5030_744889030330_33u  1  2  3  4  PARAMS:
+  Cww=21.7p
+  Rp1=21944
+  Cp1=27.563p
+  Lp1=33u
+  Rp2=183718
+  Cp2=5.313p
+  Lp2=297u
+  RDC1=1.466
+  RDC2=3.758
+  K=0.998399392428374
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
