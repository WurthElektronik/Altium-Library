**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Power Inductor
* Matchcode:              WE-PD2 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1054_744776012_1.2u 1 2
Rp 1 2 3008.47196972
Cp 1 2 1.94370161067p
Rs 1 N3 0.006
L1 N3 2 1.2u
.ends 1054_744776012_1.2u
*******
.subckt 1054_744776022_2.2u 1 2
Rp 1 2 6108.9488222
Cp 1 2 2.294256488p
Rs 1 N3 0.01
L1 N3 2 2.2u
.ends 1054_744776022_2.2u
*******
.subckt 1054_744776033_3.3u 1 2
Rp 1 2 8340.68168151
Cp 1 2 3.360864162p
Rs 1 N3 0.015
L1 N3 2 3.3u
.ends 1054_744776033_3.3u
*******
.subckt 1054_744776047_4.7u 1 2
Rp 1 2 9941.61357226
Cp 1 2 3.488313895p
Rs 1 N3 0.017
L1 N3 2 4.7u
.ends 1054_744776047_4.7u
*******
.subckt 1054_744776056_5.6u 1 2
Rp 1 2 11430.8111188
Cp 1 2 3.583689286p
Rs 1 N3 0.019
L1 N3 2 5.6u
.ends 1054_744776056_5.6u
*******
.subckt 1054_744776068_6.8u 1 2
Rp 1 2 13905.6215271
Cp 1 2 3.429901273p
Rs 1 N3 0.022
L1 N3 2 6.8u
.ends 1054_744776068_6.8u
*******
.subckt 1054_744776082_8.2u 1 2
Rp 1 2 17802.6827169
Cp 1 2 3.1792169294p
Rs 1 N3 0.026
L1 N3 2 8.2u
.ends 1054_744776082_8.2u
*******
.subckt 1054_74477610_10u 1 2
Rp 1 2 18500
Cp 1 2 3.3p
Rs 1 N3 0.0275
L1 N3 2 10u
.ends 1054_74477610_10u
*******
.subckt 1054_744776112_12u 1 2
Rp 1 2 19000
Cp 1 2 3.7p
Rs 1 N3 0.0326
L1 N3 2 12u
.ends 1054_744776112_12u
*******
.subckt 1054_744776115_15u 1 2
Rp 1 2 20000
Cp 1 2 4p
Rs 1 N3 0.034
L1 N3 2 15u
.ends 1054_744776115_15u
*******
.subckt 1054_744776118_18u 1 2
Rp 1 2 18500
Cp 1 2 4.26p
Rs 1 N3 0.0428
L1 N3 2 18u
.ends 1054_744776118_18u
*******
.subckt 1054_744776122_22u 1 2
Rp 1 2 22000
Cp 1 2 4.3p
Rs 1 N3 0.0511
L1 N3 2 22u
.ends 1054_744776122_22u
*******
.subckt 1054_744776127_27u 1 2
Rp 1 2 22000
Cp 1 2 4.7p
Rs 1 N3 0.0627
L1 N3 2 27u
.ends 1054_744776127_27u
*******
.subckt 1054_744776133_33u 1 2
Rp 1 2 28000
Cp 1 2 4.1p
Rs 1 N3 0.0826
L1 N3 2 33u
.ends 1054_744776133_33u
*******
.subckt 1054_744776139_39u 1 2
Rp 1 2 40000
Cp 1 2 4.5p
Rs 1 N3 0.0983
L1 N3 2 39u
.ends 1054_744776139_39u
*******
.subckt 1054_744776147_47u 1 2
Rp 1 2 40000
Cp 1 2 4.5p
Rs 1 N3 0.0951
L1 N3 2 47u
.ends 1054_744776147_47u
*******
.subckt 1054_744776156_56u 1 2
Rp 1 2 35000
Cp 1 2 5p
Rs 1 N3 0.112
L1 N3 2 56u
.ends 1054_744776156_56u
*******
.subckt 1054_744776168_68u 1 2
Rp 1 2 50000
Cp 1 2 5.1p
Rs 1 N3 0.138
L1 N3 2 68u
.ends 1054_744776168_68u
*******
.subckt 1054_744776182_82u 1 2
Rp 1 2 50000
Cp 1 2 5.5p
Rs 1 N3 0.15
L1 N3 2 82u
.ends 1054_744776182_82u
*******
.subckt 1054_74477620_100u 1 2
Rp 1 2 55000
Cp 1 2 5.3p
Rs 1 N3 0.2
L1 N3 2 100u
.ends 1054_74477620_100u
*******
.subckt 1054_744776212_120u 1 2
Rp 1 2 60000
Cp 1 2 5p
Rs 1 N3 0.243
L1 N3 2 120u
.ends 1054_744776212_120u
*******
.subckt 1054_744776215_150u 1 2
Rp 1 2 24000
Cp 1 2 3.59p
Rs 1 N3 0.3
L1 N3 2 150u
.ends 1054_744776215_150u
*******
.subckt 1054_744776218_180u 1 2
Rp 1 2 28700
Cp 1 2 4.13p
Rs 1 N3 0.32
L1 N3 2 180u
.ends 1054_744776218_180u
*******
.subckt 1054_744776222_220u 1 2
Rp 1 2 36000
Cp 1 2 4.72p
Rs 1 N3 0.4511
L1 N3 2 220u
.ends 1054_744776222_220u
*******
.subckt 1054_744776227_270u 1 2
Rp 1 2 85000
Cp 1 2 6.5p
Rs 1 N3 0.5
L1 N3 2 270u
.ends 1054_744776227_270u
*******
.subckt 1054_744776233_330u 1 2
Rp 1 2 110000
Cp 1 2 5.5p
Rs 1 N3 0.75
L1 N3 2 330u
.ends 1054_744776233_330u
*******
.subckt 1054_744776239_390u 1 2
Rp 1 2 120000
Cp 1 2 5.5p
Rs 1 N3 0.794
L1 N3 2 390u
.ends 1054_744776239_390u
*******
.subckt 1054_744776247_470u 1 2
Rp 1 2 150000
Cp 1 2 5.5p
Rs 1 N3 0.969
L1 N3 2 470u
.ends 1054_744776247_470u
*******
.subckt 1054_744776256_560u 1 2
Rp 1 2 170000
Cp 1 2 5.7p
Rs 1 N3 1.047
L1 N3 2 560u
.ends 1054_744776256_560u
*******
.subckt 1054_744776268_680u 1 2
Rp 1 2 190000
Cp 1 2 6.3p
Rs 1 N3 1.245
L1 N3 2 680u
.ends 1054_744776268_680u
*******
.subckt 1054_744776282_820u 1 2
Rp 1 2 210000
Cp 1 2 6.5p
Rs 1 N3 1.42
L1 N3 2 820u
.ends 1054_744776282_820u
*******
.subckt 1054_74477630_1m 1 2
Rp 1 2 226969
Cp 1 2 5.451418238p
Rs 1 N3 2.6
L1 N3 2 1000u
.ends 1054_74477630_1m
*******
.subckt 1054_744776312_1.2m 1 2
Rp 1 2 252394.564814
Cp 1 2 5.0011317632p
Rs 1 N3 3
L1 N3 2 1200u
.ends 1054_744776312_1.2m
*******
.subckt 1054_744776322_2.2m 1 2
Rp 1 2 299060.334267
Cp 1 2 6.123420137p
Rs 1 N3 5.3
L1 N3 2 2200u
.ends 1054_744776322_2.2m
*******
.subckt 3521_7447732010_1u 1 2
Rp 1 2 4178.13
Cp 1 2 1.057p
Rs 1 N3 0.039
L1 N3 2 1u
.ends 3521_7447732010_1u
*******
.subckt 3521_7447732015_1.5u 1 2
Rp 1 2 5992.2
Cp 1 2 1.004p
Rs 1 N3 0.054
L1 N3 2 1.5u
.ends 3521_7447732015_1.5u
*******
.subckt 3521_7447732022_2.2u 1 2
Rp 1 2 7841
Cp 1 2 1.016p
Rs 1 N3 0.07
L1 N3 2 2.2u
.ends 3521_7447732022_2.2u
*******
.subckt 3521_7447732033_3.3u 1 2
Rp 1 2 11393
Cp 1 2 1.133p
Rs 1 N3 0.091
L1 N3 2 3.3u
.ends 3521_7447732033_3.3u
*******
.subckt 3521_7447732047_4.7u 1 2
Rp 1 2 13076
Cp 1 2 1.104p
Rs 1 N3 0.125
L1 N3 2 4.7u
.ends 3521_7447732047_4.7u
*******
.subckt 3521_7447732068_6.8u 1 2
Rp 1 2 17163
Cp 1 2 1.368p
Rs 1 N3 0.17
L1 N3 2 6.8u
.ends 3521_7447732068_6.8u
*******
.subckt 3521_7447732110_10u 1 2
Rp 1 2 21877
Cp 1 2 1.189p
Rs 1 N3 0.237
L1 N3 2 10u
.ends 3521_7447732110_10u
*******
.subckt 3521_7447732115_15u 1 2
Rp 1 2 28826
Cp 1 2 1.334p
Rs 1 N3 0.347
L1 N3 2 15u
.ends 3521_7447732115_15u
*******
.subckt 3521_7447732122_22u 1 2
Rp 1 2 33835
Cp 1 2 1.695p
Rs 1 N3 0.561
L1 N3 2 22u
.ends 3521_7447732122_22u
*******
.subckt 3521_7447732133_33u 1 2
Rp 1 2 39684
Cp 1 2 1.749p
Rs 1 N3 0.778
L1 N3 2 33u
.ends 3521_7447732133_33u
*******
.subckt 3521_7447732147_47u 1 2
Rp 1 2 60003
Cp 1 2 1.378p
Rs 1 N3 1.11
L1 N3 2 47u
.ends 3521_7447732147_47u
*******
.subckt 3521_7447732168_68u 1 2
Rp 1 2 73284
Cp 1 2 1.492p
Rs 1 N3 1.57
L1 N3 2 68u
.ends 3521_7447732168_68u
*******
.subckt 3521_7447732210_100u 1 2
Rp 1 2 85290.4
Cp 1 2 1.41646p
Rs 1 N3 2.42
L1 N3 2 100u
.ends 3521_7447732210_100u
*******
.subckt 4532_7447730_1u 1 2
Rp 1 2 3700
Cp 1 2 1.33p
Rs 1 N3 0.014
L1 N3 2 1u
.ends 4532_7447730_1u
*******
.subckt 4532_744773014_1.4u 1 2
Rp 1 2 4550
Cp 1 2 1.83p
Rs 1 N3 0.022
L1 N3 2 1.4u
.ends 4532_744773014_1.4u
*******
.subckt 4532_744773018_1.8u 1 2
Rp 1 2 8000
Cp 1 2 2.18p
Rs 1 N3 0.028
L1 N3 2 1.8u
.ends 4532_744773018_1.8u
*******
.subckt 4532_744773022_2.2u 1 2
Rp 1 2 8750
Cp 1 2 2.5p
Rs 1 N3 0.034
L1 N3 2 2.2u
.ends 4532_744773022_2.2u
*******
.subckt 4532_744773027_2.7u 1 2
Rp 1 2 7900
Cp 1 2 1.86p
Rs 1 N3 0.039
L1 N3 2 2.7u
.ends 4532_744773027_2.7u
*******
.subckt 4532_744773033_3.3u 1 2
Rp 1 2 9800
Cp 1 2 2.16p
Rs 1 N3 0.041
L1 N3 2 3.3u
.ends 4532_744773033_3.3u
*******
.subckt 4532_744773039_3.9u 1 2
Rp 1 2 11500
Cp 1 2 1.8p
Rs 1 N3 0.054
L1 N3 2 3.9u
.ends 4532_744773039_3.9u
*******
.subckt 4532_744773047_4.7u 1 2
Rp 1 2 14200
Cp 1 2 1.95p
Rs 1 N3 0.059
L1 N3 2 4.7u
.ends 4532_744773047_4.7u
*******
.subckt 4532_744773056_5.6u 1 2
Rp 1 2 22000
Cp 1 2 1.86p
Rs 1 N3 0.069
L1 N3 2 5.6u
.ends 4532_744773056_5.6u
*******
.subckt 4532_744773068_6.8u 1 2
Rp 1 2 13300
Cp 1 2 2.14p
Rs 1 N3 0.076
L1 N3 2 6.8u
.ends 4532_744773068_6.8u
*******
.subckt 4532_744773082_8.2u 1 2
Rp 1 2 18000
Cp 1 2 2.1p
Rs 1 N3 0.116
L1 N3 2 8.2u
.ends 4532_744773082_8.2u
*******
.subckt 4532_74477310_10u 1 2
Rp 1 2 19000
Cp 1 2 2.2p
Rs 1 N3 0.118
L1 N3 2 10u
.ends 4532_74477310_10u
*******
.subckt 4532_744773112_12u 1 2
Rp 1 2 21000
Cp 1 2 2.27p
Rs 1 N3 0.156
L1 N3 2 12u
.ends 4532_744773112_12u
*******
.subckt 4532_744773115_15u 1 2
Rp 1 2 25700
Cp 1 2 2.35p
Rs 1 N3 0.204
L1 N3 2 15u
.ends 4532_744773115_15u
*******
.subckt 4532_744773118_18u 1 2
Rp 1 2 29000
Cp 1 2 2.82p
Rs 1 N3 0.225
L1 N3 2 18u
.ends 4532_744773118_18u
*******
.subckt 4532_744773122_22u 1 2
Rp 1 2 31000
Cp 1 2 2.47p
Rs 1 N3 0.261
L1 N3 2 22u
.ends 4532_744773122_22u
*******
.subckt 4532_744773127_27u 1 2
Rp 1 2 33000
Cp 1 2 2.4p
Rs 1 N3 0.328
L1 N3 2 27u
.ends 4532_744773127_27u
*******
.subckt 4532_744773133_33u 1 2
Rp 1 2 44200
Cp 1 2 2.69p
Rs 1 N3 0.37
L1 N3 2 33u
.ends 4532_744773133_33u
*******
.subckt 4532_744773139_39u 1 2
Rp 1 2 46200
Cp 1 2 2.4p
Rs 1 N3 0.418
L1 N3 2 39u
.ends 4532_744773139_39u
*******
.subckt 4532_744773147_47u 1 2
Rp 1 2 58200
Cp 1 2 2.42p
Rs 1 N3 0.523
L1 N3 2 47u
.ends 4532_744773147_47u
*******
.subckt 4532_744773156_56u 1 2
Rp 1 2 61700
Cp 1 2 2.79p
Rs 1 N3 0.714
L1 N3 2 56u
.ends 4532_744773156_56u
*******
.subckt 4532_744773168_68u 1 2
Rp 1 2 67200
Cp 1 2 2.53p
Rs 1 N3 0.754
L1 N3 2 68u
.ends 4532_744773168_68u
*******
.subckt 4532_74477330A_1000u 1 2
Rp 1 2 306000
Cp 1 2 2.334p
Rs 1 N3 1.25
L1 N3 2 1000u
.ends 4532_74477330A_1000u
*******
.subckt 5848_744774003_0.33u 1 2
Rp 1 2 1389
Cp 1 2 0.689p
Rs 1 N3 0.006
L1 N3 2 0.287u
.ends 5848_744774003_0.33u
*******
.subckt 5848_744774022_2.2u 1 2
Rp 1 2 8000
Cp 1 2 3.2p
Rs 1 N3 0.026
L1 N3 2 2.2u
.ends 5848_744774022_2.2u
*******
.subckt 5848_744774027_2.7u 1 2
Rp 1 2 10300
Cp 1 2 4.2p
Rs 1 N3 0.032
L1 N3 2 2.7u
.ends 5848_744774027_2.7u
*******
.subckt 5848_744774033_3.3u 1 2
Rp 1 2 12000
Cp 1 2 3.4p
Rs 1 N3 0.042
L1 N3 2 3.3u
.ends 5848_744774033_3.3u
*******
.subckt 5848_744774047_4.7u 1 2
Rp 1 2 14500
Cp 1 2 3.4p
Rs 1 N3 0.056
L1 N3 2 4.7u
.ends 5848_744774047_4.7u
*******
.subckt 5848_744774068_6.8u 1 2
Rp 1 2 16200
Cp 1 2 4.8p
Rs 1 N3 0.071
L1 N3 2 6.8u
.ends 5848_744774068_6.8u
*******
.subckt 5848_74477410_10u 1 2
Rp 1 2 18400
Cp 1 2 2.6p
Rs 1 N3 0.055
L1 N3 2 10u
.ends 5848_74477410_10u
*******
.subckt 5848_744774112_12u 1 2
Rp 1 2 22000
Cp 1 2 3p
Rs 1 N3 0.065
L1 N3 2 12u
.ends 5848_744774112_12u
*******
.subckt 5848_744774115_15u 1 2
Rp 1 2 29500
Cp 1 2 2.95p
Rs 1 N3 0.089
L1 N3 2 15u
.ends 5848_744774115_15u
*******
.subckt 5848_744774118_18u 1 2
Rp 1 2 31000
Cp 1 2 2.95p
Rs 1 N3 0.104
L1 N3 2 18u
.ends 5848_744774118_18u
*******
.subckt 5848_744774122_22u 1 2
Rp 1 2 26500
Cp 1 2 3.4p
Rs 1 N3 0.109
L1 N3 2 22u
.ends 5848_744774122_22u
*******
.subckt 5848_744774127_27u 1 2
Rp 1 2 35000
Cp 1 2 3.47p
Rs 1 N3 0.133
L1 N3 2 27u
.ends 5848_744774127_27u
*******
.subckt 5848_744774133_33u 1 2
Rp 1 2 38000
Cp 1 2 3.5p
Rs 1 N3 0.15
L1 N3 2 33u
.ends 5848_744774133_33u
*******
.subckt 5848_744774139_39u 1 2
Rp 1 2 45000
Cp 1 2 3.55p
Rs 1 N3 0.215
L1 N3 2 39u
.ends 5848_744774139_39u
*******
.subckt 5848_744774147_47u 1 2
Rp 1 2 52500
Cp 1 2 3.72p
Rs 1 N3 0.26
L1 N3 2 47u
.ends 5848_744774147_47u
*******
.subckt 5848_744774156_56u 1 2
Rp 1 2 53800
Cp 1 2 3.52p
Rs 1 N3 0.298
L1 N3 2 56u
.ends 5848_744774156_56u
*******
.subckt 5848_744774168_68u 1 2
Rp 1 2 54000
Cp 1 2 3.8p
Rs 1 N3 0.313
L1 N3 2 68u
.ends 5848_744774168_68u
*******
.subckt 5848_744774182_82u 1 2
Rp 1 2 66900
Cp 1 2 3.8p
Rs 1 N3 0.475
L1 N3 2 82u
.ends 5848_744774182_82u
*******
.subckt 5848_74477420_100u 1 2
Rp 1 2 95000
Cp 1 2 3.89p
Rs 1 N3 0.51
L1 N3 2 100u
.ends 5848_74477420_100u
*******
.subckt 5848_744774212_120u 1 2
Rp 1 2 89000
Cp 1 2 3.7p
Rs 1 N3 0.66
L1 N3 2 120u
.ends 5848_744774212_120u
*******
.subckt 5848_744774215_150u 1 2
Rp 1 2 90500
Cp 1 2 3.8p
Rs 1 N3 0.72
L1 N3 2 150u
.ends 5848_744774215_150u
*******
.subckt 5848_744774218_180u 1 2
Rp 1 2 105000
Cp 1 2 4.1p
Rs 1 N3 0.85
L1 N3 2 180u
.ends 5848_744774218_180u
*******
.subckt 5848_744774222_220u 1 2
Rp 1 2 110000
Cp 1 2 4.2p
Rs 1 N3 0.945
L1 N3 2 220u
.ends 5848_744774222_220u
*******
.subckt 7850_744775022_2.2u 1 2
Rp 1 2 5872.78138167
Cp 1 2 2.65935962351p
Rs 1 N3 0.015
L1 N3 2 2.2u
.ends 7850_744775022_2.2u
*******
.subckt 7850_744775033_3.3u 1 2
Rp 1 2 8518.85993879
Cp 1 2 2.7034855228p
Rs 1 N3 0.018
L1 N3 2 3.3u
.ends 7850_744775033_3.3u
*******
.subckt 7850_744775047_4.7u 1 2
Rp 1 2 11042.0212798
Cp 1 2 3.46979460166p
Rs 1 N3 0.019
L1 N3 2 4.7u
.ends 7850_744775047_4.7u
*******
.subckt 7850_744775056_5.6u 1 2
Rp 1 2 12712.0393799
Cp 1 2 3.26388455702p
Rs 1 N3 0.022
L1 N3 2 5.6u
.ends 7850_744775056_5.6u
*******
.subckt 7850_744775068_6.8u 1 2
Rp 1 2 13285.326443
Cp 1 2 3.58505630156p
Rs 1 N3 0.026
L1 N3 2 6.8u
.ends 7850_744775068_6.8u
*******
.subckt 7850_744775082_8.2u 1 2
Rp 1 2 16359.5409893
Cp 1 2 3.46552296283p
Rs 1 N3 0.04
L1 N3 2 8.2u
.ends 7850_744775082_8.2u
*******
.subckt 7850_74477510_10u 1 2
Rp 1 2 15000
Cp 1 2 3p
Rs 1 N3 0.04
L1 N3 2 10u
.ends 7850_74477510_10u
*******
.subckt 7850_744775112_12u 1 2
Rp 1 2 29000
Cp 1 2 4.02p
Rs 1 N3 0.0417
L1 N3 2 12u
.ends 7850_744775112_12u
*******
.subckt 7850_744775115_15u 1 2
Rp 1 2 19000
Cp 1 2 3.86p
Rs 1 N3 0.0439
L1 N3 2 15u
.ends 7850_744775115_15u
*******
.subckt 7850_744775118_18u 1 2
Rp 1 2 21000
Cp 1 2 3.7p
Rs 1 N3 0.0526
L1 N3 2 18u
.ends 7850_744775118_18u
*******
.subckt 7850_744775122_22u 1 2
Rp 1 2 21000
Cp 1 2 4p
Rs 1 N3 0.0654
L1 N3 2 22u
.ends 7850_744775122_22u
*******
.subckt 7850_744775127_27u 1 2
Rp 1 2 25000
Cp 1 2 3.4p
Rs 1 N3 0.0738
L1 N3 2 27u
.ends 7850_744775127_27u
*******
.subckt 7850_744775133_33u 1 2
Rp 1 2 30000
Cp 1 2 4.7p
Rs 1 N3 0.0878
L1 N3 2 33u
.ends 7850_744775133_33u
*******
.subckt 7850_744775139_39u 1 2
Rp 1 2 35000
Cp 1 2 4.8p
Rs 1 N3 0.116
L1 N3 2 39u
.ends 7850_744775139_39u
*******
.subckt 7850_744775147_47u 1 2
Rp 1 2 40000
Cp 1 2 4p
Rs 1 N3 0.1343
L1 N3 2 47u
.ends 7850_744775147_47u
*******
.subckt 7850_744775156_56u 1 2
Rp 1 2 35000
Cp 1 2 4.55p
Rs 1 N3 0.189
L1 N3 2 56u
.ends 7850_744775156_56u
*******
.subckt 7850_744775168_68u 1 2
Rp 1 2 55000
Cp 1 2 3.8p
Rs 1 N3 0.218
L1 N3 2 68u
.ends 7850_744775168_68u
*******
.subckt 7850_744775182_82u 1 2
Rp 1 2 60000
Cp 1 2 4.25p
Rs 1 N3 0.208
L1 N3 2 82u
.ends 7850_744775182_82u
*******
.subckt 7850_74477520_100u 1 2
Rp 1 2 65000
Cp 1 2 4.3p
Rs 1 N3 0.2482
L1 N3 2 100u
.ends 7850_74477520_100u
*******
.subckt 7850_744775210_120u 1 2
Rp 1 2 58000
Cp 1 2 4.5p
Rs 1 N3 0.308
L1 N3 2 120u
.ends 7850_744775210_120u
*******
.subckt 7850_744775215_150u 1 2
Rp 1 2 95000
Cp 1 2 4.2p
Rs 1 N3 0.4666
L1 N3 2 150u
.ends 7850_744775215_150u
*******
.subckt 7850_744775218_180u 1 2
Rp 1 2 105000
Cp 1 2 4.5p
Rs 1 N3 0.5741
L1 N3 2 180u
.ends 7850_744775218_180u
*******
.subckt 7850_744775222_220u 1 2
Rp 1 2 95000
Cp 1 2 4.4p
Rs 1 N3 0.614
L1 N3 2 220u
.ends 7850_744775222_220u
*******
.subckt 7850_744775227_270u 1 2
Rp 1 2 100000
Cp 1 2 5p
Rs 1 N3 0.699
L1 N3 2 270u
.ends 7850_744775227_270u
*******
.subckt 7850_744775233_330u 1 2
Rp 1 2 110000
Cp 1 2 5.3p
Rs 1 N3 0.81
L1 N3 2 330u
.ends 7850_744775233_330u
*******
.subckt 7850_744775239_390u 1 2
Rp 1 2 180000
Cp 1 2 5p
Rs 1 N3 1.151
L1 N3 2 390u
.ends 7850_744775239_390u
*******
.subckt 7850_744775247_470u 1 2
Rp 1 2 165000
Cp 1 2 5p
Rs 1 N3 1.37
L1 N3 2 470u
.ends 7850_744775247_470u
*******
.subckt 7850_74477530_1m 1 2
Rp 1 2 187304.915771
Cp 1 2 4.36976277949p
Rs 1 N3 3.3
L1 N3 2 1000u
.ends 7850_74477530_1m
*******
.subckt 1054_744776260_600u 1 2
Rp 1 2 180000
Cp 1 2 5p
Rs 1 N3 1
L1 N3 2 570u
.ends 1054_744776260_600u