**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Multilayer Ceramic SMT Inductor
* Matchcode:              WE-MCI
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-23
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0402_7847803100_1n 1 2
C1 1 N7 250.4375f
L1 1 N1 0.95n
L2 N1 N2 67.3802p
L3 N2 N3 322.6669p
L4 N3 N4 451.7293p
L5 N4 N5 77.2222p
L6 N5 N6 54.4474p
R1 2 N1 325.1654m
R2 2 N2 150.2242m
R3 2 N3 424.1842m
R4 2 N4 391.6119m
R5 2 N5 348.2740m
R6 2 N6 96.5700m
R7 2 N7 1.9664
R8 2 1 10g
.ends 
*******
.subckt 0402_7847803270_2.7n 1 2
C1 1 N7 328.2021f
L1 1 N1 2.55n
L2 N1 N2 211.0089p
L3 N2 N3 308.5137p
L4 N3 N4 434.6384p
L5 N4 N5 77.1557p
L6 N5 N6 54.4297p
R1 2 N1 512.1942m
R2 2 N2 279.7939m
R3 2 N3 409.8297m
R4 2 N4 396.9486m
R5 2 N5 356.5497m
R6 2 N6 97.6827m
R7 2 N7 1.9689
R8 2 1 10g
.ends 
*******
.subckt 0402_7847803330_3.3n 1 2
C1 1 N7 279.6563f
L1 1 N1 3.1n
L2 N1 N2 195.7892p
L3 N2 N3 548.9631p
L4 N3 N4 709.8211p
L5 N4 N5 79.2776p
L6 N5 N6 55.8162p
R1 2 N1 806.2502m
R2 2 N2 451.7123m
R3 2 N3 525.1138m
R4 2 N4 531.1421m
R5 2 N5 502.9249m
R6 2 N6 118.1228m
R7 2 N7 1.9691
R8 2 1 10g
.ends 
*******
.subckt 0402_7847803390_3.9n 1 2
C1 1 N7 402.3598f
L1 1 N1 3.72n
L2 N1 N2 331.8377p
L3 N2 N3 649.2075p
L4 N3 N4 823.1100p
L5 N4 N5 80.1764p
L6 N5 N6 56.4343p
R1 2 N1 809.8159m
R2 2 N2 627.9723m
R3 2 N3 574.3743m
R4 2 N4 592.1578m
R5 2 N5 566.4181m
R6 2 N6 129.2745m
R7 2 N7 1.9722
R8 2 1 10g
.ends 
*******
.subckt 0402_7847803560_5.6n 1 2
C1 1 N7 383.7784f
L1 1 N1 5.3n
L2 N1 N2 593.7969p
L3 N2 N3 784.7160p
L4 N3 N4 985.5525p
L5 N4 N5 81.4082p
L6 N5 N6 57.2765p
R1 2 N1 1.0909
R2 2 N2 627.3629m
R3 2 N3 671.9811m
R4 2 N4 661.5756m
R5 2 N5 636.2967m
R6 2 N6 142.2376m
R7 2 N7 1.9698
R8 2 1 10g
.ends 
*******
.subckt 0402_7847803680_6.8n 1 2
C1 1 N7 291.8149f
L1 1 N1 6.5n
L2 N1 N2 723.5885p
L3 N2 N3 1.1901n
L4 N3 N4 1.3769n
L5 N4 N5 84.3277p
L6 N5 N6 59.2644p
R1 2 N1 1.2076
R2 2 N2 728.6026m
R3 2 N3 944.0779m
R4 2 N4 838.8510m
R5 2 N5 814.8120m
R6 2 N6 176.7420m
R7 2 N7 1.9647
R8 2 1 10g
.ends 
*******
.subckt 0402_7847803820_8.2n 1 2
C1 1 N7 283.9689f
L1 1 N1 7.7n
L2 N1 N2 924.9233p
L3 N2 N3 1.6741n
L4 N3 N4 1.8632n
L5 N4 N5 87.9572p
L6 N5 N6 61.7488p
R1 2 N1 1.8774
R2 2 N2 867.0091m
R3 2 N3 1.2342
R4 2 N4 1.08
R5 2 N5 1.0575
R6 2 N6 226.9601m
R7 2 N7 2.9576
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804100_10n 1 2
C1 1 N7 283.9689f
L1 1 N1 9.3n
L2 N1 N2 1.0519n
L3 N2 N3 1.9021n
L4 N3 N4 2.0582n
L5 N4 N5 87.9880p
L6 N5 N6 61.7821p
R1 2 N1 1.9992
R2 2 N2 891.6052m
R3 2 N3 1.2352
R4 2 N4 1.0817
R5 2 N5 1.0592
R6 2 N6 262.2584m
R7 2 N7 2.9628
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804101_100n 1 2
C1 1 N7 230.2332f
L1 1 N1 90n
L2 N1 N2 9.5700n
L3 N2 N3 19.2563n
L4 N3 N4 20.8626n
L5 N4 N5 92.6028p
L6 N5 N6 65.4207p
R1 2 N1 21.3883
R2 2 N2 7.1149
R3 2 N3 4.3109
R4 2 N4 2.9427
R5 2 N5 2.9357
R6 2 N6 2.5456
R7 2 N7 5.6084
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804120_12n 1 2
C1 1 N7 194.5952f
L1 1 N1 11n
L2 N1 N2 1.3585n
L3 N2 N3 3.0908n
L4 N3 N4 3.2821n
L5 N4 N5 91.5040p
L6 N5 N6 64.7058p
R1 2 N1 2.8113
R2 2 N2 904.4775m
R3 2 N3 1.2507
R4 2 N4 1.0999
R5 2 N5 1.0778
R6 2 N6 437.2241m
R7 2 N7 2.9866
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804150_15n 1 2
C1 1 N7 207.3289f
L1 1 N1 13.5n
L2 N1 N2 1.7941n
L3 N2 N3 4.5924n
L4 N3 N4 4.1124n
L5 N4 N5 91.5584p
L6 N5 N6 64.7365p
R1 2 N1 3.4834
R2 2 N2 997.4626m
R3 2 N3 1.2709
R4 2 N4 1.1133
R5 2 N5 1.0916
R6 2 N6 511.9220m
R7 2 N7 3.0122
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804180_18n 1 2
C1 1 N7 202.5706f
L1 1 N1 16.5n
L2 N1 N2 1.9675n
L3 N2 N3 5.0093n
L4 N3 N4 5.1131n
L5 N4 N5 91.6163p
L6 N5 N6 64.7606p
R1 2 N1 3.9793
R2 2 N2 1.505
R3 2 N3 1.2899
R4 2 N4 1.1703
R5 2 N5 1.1505
R6 2 N6 724.0214m
R7 2 N7 3.1349
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804181_180n 1 2
C1 1 N7 323.1487f
L1 1 N1 160n
L2 N1 N2 23.0017n
L3 N2 N3 49.1098n
L4 N3 N4 207.9221n
L5 N4 N5 94.0227p
L6 N5 N6 67.2068p
R1 2 N1 27.3466
R2 2 N2 9.8039
R3 2 N3 4.1216
R4 2 N4 3.3756
R5 2 N5 3.3698
R6 2 N6 3.0907
R7 2 N7 6.3753
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804270_27n 1 2
C1 1 N7 176.5554f
L1 1 N1 25n
L2 N1 N2 3.4691n
L3 N2 N3 8.3863n
L4 N3 N4 10.8230n
L5 N4 N5 91.7217p
L6 N5 N6 64.5940p
R1 2 N1 6.6329
R2 2 N2 2.3043
R3 2 N3 1.5061
R4 2 N4 1.4488
R5 2 N5 1.4349
R6 2 N6 1.2342
R7 2 N7 3.6389
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804271_270n 1 2
C1 1 N7 474.3076f
L1 1 N1 230n
L2 N1 N2 49.4235n
L3 N2 N3 189.2132n
L4 N3 N4 207.9221n
L5 N4 N5 92.9865p
L6 N5 N6 65.2852p
R1 2 N1 28.9698
R2 2 N2 7.8952
R3 2 N3 5.8641
R4 2 N4 4.009
R5 2 N5 4.0042
R6 2 N6 3.8288
R7 2 N7 16.4566
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804330_33n 1 2
C1 1 N7 180.6446f
L1 1 N1 31n
L2 N1 N2 4.3162n
L3 N2 N3 8.5019n
L4 N3 N4 10.9030n
L5 N4 N5 91.7258p
L6 N5 N6 64.5955p
R1 2 N1 6.6824
R2 2 N2 2.3107
R3 2 N3 1.5114
R4 2 N4 1.4523
R5 2 N5 1.4384
R6 2 N6 1.239
R7 2 N7 3.6611
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804390_39n 1 2
C1 1 N7 179.9775f
L1 1 N1 36.5n
L2 N1 N2 5.2312n
L3 N2 N3 13.5132n
L4 N3 N4 14.7242n
L5 N4 N5 91.7075p
L6 N5 N6 64.3636p
R1 2 N1 8.3342
R2 2 N2 2.6616
R3 2 N3 1.7671
R4 2 N4 1.6359
R5 2 N5 1.6242
R6 2 N6 1.4787
R7 2 N7 4.0193
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804470_47n 1 2
C1 1 N7 210.5192f
L1 1 N1 43n
L2 N1 N2 5.0495n
L3 N2 N3 9.4856n
L4 N3 N4 20.3991n
L5 N4 N5 92.3790p
L6 N5 N6 64.8352p
R1 2 N1 9.4594
R2 2 N2 4.1477
R3 2 N3 2.1457
R4 2 N4 2.3175
R5 2 N5 2.3108
R6 2 N6 2.2515
R7 2 N7 9.2499
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804560_56n 1 2
C1 1 N7 240.5192f
L1 1 N1 52n
L2 N1 N2 7.0551n
L3 N2 N3 12.5903n
L4 N3 N4 20.3991n
L5 N4 N5 92.6307p
L6 N5 N6 64.9042p
R1 2 N1 10.5992
R2 2 N2 4.0413
R3 2 N3 2.6169
R4 2 N4 2.5454
R5 2 N5 2.5391
R6 2 N6 2.4907
R7 2 N7 9.4944
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804680_68n 1 2
C1 1 N7 228.9714f
L1 1 N1 63n
L2 N1 N2 8.5654n
L3 N2 N3 15.2978n
L4 N3 N4 20.3991n
L5 N4 N5 93.3419p
L6 N5 N6 65.6314p
R1 2 N1 11.3757
R2 2 N2 3.9293
R3 2 N3 2.9744
R4 2 N4 2.8492
R5 2 N5 2.8435
R6 2 N6 2.6137
R7 2 N7 9.8426
R8 2 1 10g
.ends 
*******
.subckt 0402_7847804820_82n 1 2
C1 1 N7 290.9087f
L1 1 N1 76n
L2 N1 N2 10.3090n
L3 N2 N3 18.6637n
L4 N3 N4 20.3991n
L5 N4 N5 96.9908p
L6 N5 N6 68.3809p
R1 2 N1 14.2916
R2 2 N2 5.5482
R3 2 N3 4.8936
R4 2 N4 4.431
R5 2 N5 4.4251
R6 2 N6 2.6137
R7 2 N7 9.969
R8 2 1 10g
.ends 
*******
.subckt 0603_7847805100_1n 1 2
C1 1 N7 286.0060f
L1 1 N1 0.95n
L2 N1 N2 36.3973p
L3 N2 N3 110.3289p
L4 N3 N4 322.6993p
L5 N4 N5 76.5477p
L6 N5 N6 54.0923p
R1 2 N1 165.9532m
R2 2 N2 70.5967m
R3 2 N3 216.8744m
R4 2 N4 376.1808m
R5 2 N5 340.0279m
R6 2 N6 96.0037m
R7 2 N7 1.9858
R8 2 1 10g
.ends 
*******
.subckt 0603_7847805220_2.2n 1 2
C1 1 N7 686.0925f
L1 1 N1 2.1n
L2 N1 N2 136.0516p
L3 N2 N3 166.0962p
L4 N3 N4 524.5172p
L5 N4 N5 77.7100p
L6 N5 N6 54.7805p
R1 2 N1 276.0085m
R2 2 N2 184.4143m
R3 2 N3 115.4778m
R4 2 N4 391.2767m
R5 2 N5 342.0058m
R6 2 N6 95.2030m
R7 2 N7 2.0158
R8 2 1 10g
.ends 
*******
.subckt 0603_7847805390_3.9n 1 2
C1 1 N7 398.0912f
L1 1 N1 3.8n
L2 N1 N2 182.6841p
L3 N2 N3 193.5080p
L4 N3 N4 578.7244p
L5 N4 N5 78.0710p
L6 N5 N6 55.0703p
R1 2 N1 372.9908m
R2 2 N2 228.4273m
R3 2 N3 133.9181m
R4 2 N4 404.7694m
R5 2 N5 354.5175m
R6 2 N6 96.3931m
R7 2 N7 2.0226
R8 2 1 10g
.ends 
*******
.subckt 0603_7847805470_4.7n 1 2
C1 1 N7 203.9559f
L1 1 N1 4.5n
L2 N1 N2 138.5648p
L3 N2 N3 481.1173p
L4 N3 N4 1.8998n
L5 N4 N5 85.0038p
L6 N5 N6 59.4273p
R1 2 N1 1.2702
R2 2 N2 535.5083m
R3 2 N3 417.6056m
R4 2 N4 661.5905m
R5 2 N5 613.1207m
R6 2 N6 257.2973m
R7 2 N7 3.5339
R8 2 1 10g
.ends 
*******
.subckt 0603_7847805560_5.6n 1 2
C1 1 N7 262.2938f
L1 1 N1 5.4n
L2 N1 N2 179.6066p
L3 N2 N3 482.3239p
L4 N3 N4 1.8475n
L5 N4 N5 85.0007p
L6 N5 N6 59.4256p
R1 2 N1 1.275
R2 2 N2 543.1002m
R3 2 N3 412.7223m
R4 2 N4 661.5712m
R5 2 N5 613.1259m
R6 2 N6 257.4006m
R7 2 N7 3.5349
R8 2 1 10g
.ends 
*******
.subckt 0603_7847805680_6.8n 1 2
C1 1 N7 187.3994f
L1 1 N1 6.6n
L2 N1 N2 154.5973p
L3 N2 N3 622.5872p
L4 N3 N4 2.0356n
L5 N4 N5 85.0209p
L6 N5 N6 59.4462p
R1 2 N1 1.3122
R2 2 N2 808.2573m
R3 2 N3 468.4338m
R4 2 N4 660.6548m
R5 2 N5 611.9458m
R6 2 N6 249.7392m
R7 2 N7 3.5337
R8 2 1 10g
.ends 
*******
.subckt 0603_7847805820_8.2n 1 2
C1 1 N7 263.4651f
L1 1 N1 7.9n
L2 N1 N2 413.2566p
L3 N2 N3 578.9545p
L4 N3 N4 2.3988n
L5 N4 N5 85.0380p
L6 N5 N6 59.4515p
R1 2 N1 1.372
R2 2 N2 694.2462m
R3 2 N3 505.7731m
R4 2 N4 659.6326m
R5 2 N5 610.5638m
R6 2 N6 240.6432m
R7 2 N7 3.5365
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806100_10n 1 2
C1 1 N7 305.1360f
L1 1 N1 9.5n
L2 N1 N2 503.0163p
L3 N2 N3 736.4737p
L4 N3 N4 3.5021n
L5 N4 N5 85.1487p
L6 N5 N6 59.5474p
R1 2 N1 1.5593
R2 2 N2 835.1170m
R3 2 N3 677.0231m
R4 2 N4 685.9364m
R5 2 N5 640.4659m
R6 2 N6 379.1923m
R7 2 N7 3.572
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806101_100n 1 2
C1 1 N7 304.1344f
L1 1 N1 90n
L2 N1 N2 8.1272n
L3 N2 N3 11.1356n
L4 N3 N4 23.6461n
L5 N4 N5 92.9091p
L6 N5 N6 68.1992p
R1 2 N1 10.2781
R2 2 N2 4.1769
R3 2 N3 3.283
R4 2 N4 3.6787
R5 2 N5 3.6749
R6 2 N6 1.5878
R7 2 N7 4.6827
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806120_12n 1 2
C1 1 N7 253.6627f
L1 1 N1 11.2n
L2 N1 N2 668.0841p
L3 N2 N3 755.6386p
L4 N3 N4 3.4318n
L5 N4 N5 85.1493p
L6 N5 N6 59.5524p
R1 2 N1 1.6003
R2 2 N2 888.1752m
R3 2 N3 679.1046m
R4 2 N4 686.4507m
R5 2 N5 641.0902m
R6 2 N6 380.9428m
R7 2 N7 3.5722
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806121_120n 1 2
C1 1 N7 294.1902f
L1 1 N1 105n
L2 N1 N2 9.8967n
L3 N2 N3 13.3819n
L4 N3 N4 32.6578n
L5 N4 N5 96.5566p
L6 N5 N6 73.1552p
R1 2 N1 12.5156
R2 2 N2 4.0854
R3 2 N3 3.1405
R4 2 N4 3.912
R5 2 N5 3.9087
R6 2 N6 2.4905
R7 2 N7 6.3033
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806150_15n 1 2
C1 1 N7 287.6045f
L1 1 N1 14.2n
L2 N1 N2 795.0234p
L3 N2 N3 935.0650p
L4 N3 N4 3.2890n
L5 N4 N5 85.2238p
L6 N5 N6 59.6668p
R1 2 N1 2.0627
R2 2 N2 1.0609
R3 2 N3 730.0407m
R4 2 N4 720.6483m
R5 2 N5 679.9529m
R6 2 N6 475.3827m
R7 2 N7 3.7856
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806151_150n 1 2
C1 1 N7 294.1902f
L1 1 N1 135n
L2 N1 N2 13.8160n
L3 N2 N3 14.6031n
L4 N3 N4 43.8459n
L5 N4 N5 96.5772p
L6 N5 N6 73.1769p
R1 2 N1 12.5182
R2 2 N2 4.1674
R3 2 N3 3.1726
R4 2 N4 3.9146
R5 2 N5 3.9112
R6 2 N6 2.4967
R7 2 N7 6.3052
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806180_18n 1 2
C1 1 N7 251.2455f
L1 1 N1 17.2n
L2 N1 N2 1.2044n
L3 N2 N3 1.0011n
L4 N3 N4 3.7512n
L5 N4 N5 85.2573p
L6 N5 N6 59.6897p
R1 2 N1 2.2197
R2 2 N2 1.1982
R3 2 N3 780.7182m
R4 2 N4 726.0058m
R5 2 N5 685.7112m
R6 2 N6 486.7801m
R7 2 N7 3.7885
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806181_180n 1 2
C1 1 N7 331.6229f
L1 1 N1 165n
L2 N1 N2 16.7049n
L3 N2 N3 29.9436n
L4 N3 N4 45.1320n
L5 N4 N5 91.7470p
L6 N5 N6 66.7609p
R1 2 N1 15.4465
R2 2 N2 4.7757
R3 2 N3 3.6488
R4 2 N4 4.0392
R5 2 N5 4.036
R6 2 N6 2.7987
R7 2 N7 7.0614
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806220_22n 1 2
C1 1 N7 268.7211f
L1 1 N1 21n
L2 N1 N2 1.8749n
L3 N2 N3 1.1989n
L4 N3 N4 8.3851n
L5 N4 N5 85.6932p
L6 N5 N6 60.0576p
R1 2 N1 3.0798
R2 2 N2 1.465
R3 2 N3 1.1252
R4 2 N4 812.3870m
R5 2 N5 779.3150m
R6 2 N6 654.5361m
R7 2 N7 3.8597
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806221_220n 1 2
C1 1 N7 358.9992f
L1 1 N1 200n
L2 N1 N2 21.3193n
L3 N2 N3 30.9336n
L4 N3 N4 48.6997n
L5 N4 N5 82.1985p
L6 N5 N6 53.2169p
R1 2 N1 18.9514
R2 2 N2 6.6007
R3 2 N3 5.292
R4 2 N4 4.5161
R5 2 N5 4.513
R6 2 N6 3.7845
R7 2 N7 8.0867
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806270_27n 1 2
C1 1 N7 305.5461f
L1 1 N1 25.7n
L2 N1 N2 1.9258n
L3 N2 N3 1.4003n
L4 N3 N4 8.1704n
L5 N4 N5 86.0132p
L6 N5 N6 60.5280p
R1 2 N1 3.3256
R2 2 N2 1.7003
R3 2 N3 1.3535
R4 2 N4 901.9617m
R5 2 N5 875.6226m
R6 2 N6 783.0071m
R7 2 N7 4.1152
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806271_270n 1 2
C1 1 N7 385.8094f
L1 1 N1 250n
L2 N1 N2 28.8797n
L3 N2 N3 52.9905n
L4 N3 N4 95.0048n
L5 N4 N5 82.3383p
L6 N5 N6 53.4052p
R1 2 N1 21.9132
R2 2 N2 6.817
R3 2 N3 5.2934
R4 2 N4 4.5872
R5 2 N5 4.5774
R6 2 N6 3.8751
R7 2 N7 8.131
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806330_33n 1 2
C1 1 N7 370.3324f
L1 1 N1 31.5n
L2 N1 N2 2.6951n
L3 N2 N3 1.5576n
L4 N3 N4 9.2709n
L5 N4 N5 86.0925p
L6 N5 N6 60.5822p
R1 2 N1 3.8537
R2 2 N2 2.0098
R3 2 N3 1.5207
R4 2 N4 954.7682m
R5 2 N5 931.0453m
R6 2 N6 851.3184m
R7 2 N7 4.1609
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806331_330n 1 2
C1 1 N7 384.0164f
L1 1 N1 300n
L2 N1 N2 29.2864n
L3 N2 N3 53.1097n
L4 N3 N4 147.1375n
L5 N4 N5 82.5828p
L6 N5 N6 53.7756p
R1 2 N1 25.5914
R2 2 N2 6.8479
R3 2 N3 5.2745
R4 2 N4 4.6053
R5 2 N5 4.5953
R6 2 N6 3.9073
R7 2 N7 8.1721
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806390_39n 1 2
C1 1 N7 280.2523f
L1 1 N1 37n
L2 N1 N2 3.0578n
L3 N2 N3 1.5908n
L4 N3 N4 9.9232n
L5 N4 N5 91.1086p
L6 N5 N6 67.5536p
R1 2 N1 4.6382
R2 2 N2 2.4362
R3 2 N3 2.3004
R4 2 N4 1.7454
R5 2 N5 1.7414
R6 2 N6 1.4878
R7 2 N7 2.2001
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806391_390n 1 2
C1 1 N7 366.4287f
L1 1 N1 370n
L2 N1 N2 37.0626n
L3 N2 N3 74.2171n
L4 N3 N4 446.3201n
L5 N4 N5 82.6238p
L6 N5 N6 53.8367p
R1 2 N1 25.1442
R2 2 N2 7.622
R3 2 N3 4.9299
R4 2 N4 4.6177
R5 2 N5 4.6077
R6 2 N6 3.9245
R7 2 N7 18.3647
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806470_47n 1 2
C1 1 N7 265.7943f
L1 1 N1 44n
L2 N1 N2 3.4470n
L3 N2 N3 2.2886n
L4 N3 N4 10.9051n
L5 N4 N5 90.3825p
L6 N5 N6 66.5197p
R1 2 N1 6.251
R2 2 N2 3.5406
R3 2 N3 2.9239
R4 2 N4 1.9556
R5 2 N5 1.9522
R6 2 N6 1.4878
R7 2 N7 3.0825
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806471_470n 1 2
C1 1 N7 471.9161f
L1 1 N1 435n
L2 N1 N2 55.1192n
L3 N2 N3 105.0695n
L4 N3 N4 444.4273n
L5 N4 N5 82.7210p
L6 N5 N6 53.9859p
R1 2 N1 25.6732
R2 2 N2 7.7167
R3 2 N3 4.8823
R4 2 N4 4.6197
R5 2 N5 4.6097
R6 2 N6 3.9272
R7 2 N7 18.3946
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806560_56n 1 2
C1 1 N7 313.2175f
L1 1 N1 52n
L2 N1 N2 4.4103n
L3 N2 N3 2.4209n
L4 N3 N4 11.8782n
L5 N4 N5 90.4285p
L6 N5 N6 66.5326p
R1 2 N1 6.9851
R2 2 N2 3.793
R3 2 N3 2.9239
R4 2 N4 1.9727
R5 2 N5 1.9692
R6 2 N6 1.4878
R7 2 N7 3.3285
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806680_68n 1 2
C1 1 N7 260.5880f
L1 1 N1 64n
L2 N1 N2 4.4103n
L3 N2 N3 3.2006n
L4 N3 N4 16.0855n
L5 N4 N5 92.9466p
L6 N5 N6 68.2563p
R1 2 N1 8.4935
R2 2 N2 4.1192
R3 2 N3 2.9239
R4 2 N4 3.6364
R5 2 N5 3.6325
R6 2 N6 1.2754
R7 2 N7 4.2239
R8 2 1 10g
.ends 
*******
.subckt 0603_7847806820_82n 1 2
C1 1 N7 319.6008f
L1 1 N1 77n
L2 N1 N2 7.5542n
L3 N2 N3 4.1678n
L4 N3 N4 21.6188n
L5 N4 N5 92.9485p
L6 N5 N6 68.2560p
R1 2 N1 8.5042
R2 2 N2 4.1365
R3 2 N3 2.9358
R4 2 N4 3.6367
R5 2 N5 3.6328
R6 2 N6 1.278
R7 2 N7 4.2253
R8 2 1 10g
.ends 
*******
