**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 THT High Current Inductor 
* Matchcode:             WE-HIDA
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/9/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1480_7444011480082_8.2u 1 2
Rp 1 2 3751.4
Cp 1 2 7.5266p
Rs 1 N3 0.009
L1 N3 2 7.6456u
.ends 1480_7444011480082_8.2u
*******
.subckt 1480_7444011480100_10u 1 2
Rp 1 2 3786.6
Cp 1 2 7.4402p
Rs 1 N3 0.009
L1 N3 2 8.7606u
.ends 1480_7444011480100_10u
*******
.subckt 1480_7444011480150_15u 1 2
Rp 1 2 4848.2
Cp 1 2 10.2028p
Rs 1 N3 0.01
L1 N3 2 13.7286u
.ends 1480_7444011480150_15u
*******
.subckt 1480_7444011480220_22u 1 2
Rp 1 2 5250.6
Cp 1 2 11.2868p
Rs 1 N3 0.01
L1 N3 2 20.6298u
.ends 1480_7444011480220_22u
*******
.subckt 1715_7444011715220_22u 1 2
Rp 1 2 4884.6
Cp 1 2 7.5382p
Rs 1 N3 0.007
L1 N3 2 20.7846u
.ends 1715_7444011715220_22u
*******
.subckt 1715_7444011715150_15u 1 2
Rp 1 2 4503.2
Cp 1 2 8.0702p
Rs 1 N3 0.007
L1 N3 2 14.606u
.ends 1715_7444011715150_15u
*******
.subckt 1715_7444011715100_10u 1 2
Rp 1 2 4101.6
Cp 1 2 6.582p
Rs 1 N3 0.007
L1 N3 2 8.52u
.ends 1715_7444011715100_10u
*******
.subckt 1715_7444011715082_8.2u 1 2
Rp 1 2 3901.2
Cp 1 2 7.8626p
Rs 1 N3 0.007
L1 N3 2 6.9308u
.ends 1715_7444011715082_8.2u
*******
.subckt 3119_7444013119082_8.2u 1 2
Rp 1 2 1000
Cp 1 2 11.2p
Rs 1 N3 0.0025
L1 N3 2 7.6u
.ends 3119_7444013119082_8.2u
*******
.subckt 3119_7444013119100_10u 1 2
Rp 1 2 4000
Cp 1 2 13.6666666666667p
Rs 1 N3 0.0048
L1 N3 2 10u
.ends 3119_7444013119100_10u
*******
.subckt 3119_7444013119220_22u 1 2
Rp 1 2 5000
Cp 1 2 12p
Rs 1 N3 0.0053
L1 N3 2 20u
.ends 3119_7444013119220_22u
*******
.subckt 3119_7444013119150_15u 1 2
Rp 1 2 4000
Cp 1 2 13p
Rs 1 N3 0.0048
L1 N3 2 14u
.ends 3119_7444013119150_15u
*******
.subckt 1415_7444211415082_8.2u 1 2 3 4
L1 1 N1 7.433u
Rdc1 N1 4 9.2m
Cp1 1 4 8.399p
Rp1 1 4 2314
L2 2 N2 7.433u
Rdc2  N2 3 9.2m
Cp2 2 3 8.399p
Rp2 2 3 2314
Rg1 1 0 500meg
Rg2 2 0 500meg
Rg3 3 0 500meg
Rg4 4 0 500meg
.ends
*******
.subckt 1415_7444211415100_10u 1 2 3 4
L1 1 N1 9.038u
Rdc1 N1 4 9.2m
Cp1 1 4 9.155p
Rp1 1 4 2396
L2 2 N2 9.038u
Rdc2  N2 3 9.2m
Cp2 2 3 9.155p
Rp2 2 3 2396
Rg1 1 0 500meg
Rg2 2 0 500meg
Rg3 3 0 500meg
Rg4 4 0 500meg
.ends
*******
.subckt 1415_7444211415150_15u 1 2 3 4
L1 1 N1 13.628u
Rdc1 N1 4 14.6m
Cp1 1 4 11.718p
Rp1 1 4 2908
L2 2 N2 13.628u
Rdc2  N2 3 14.6m
Cp2 2 3 11.718p
Rp2 2 3 2908
Rg1 1 0 500meg
Rg2 2 0 500meg
Rg3 3 0 500meg
Rg4 4 0 500meg
.ends
*******
.subckt 1415_7444211415220_22u 1 2 3 4
L1 1 N1 19.457u
Rdc1 N1 4 14.8m
Cp1 1 4 11.402p
Rp1 1 4 3381
L2 2 N2 19.457u
Rdc2  N2 3 14.8m
Cp2 2 3 11.402p
Rp2 2 3 3381
Rg1 1 0 500meg
Rg2 2 0 500meg
Rg3 3 0 500meg
Rg4 4 0 500meg
.ends
*******
.subckt 1521_74441521082_8.2u 1 2 3 4
L1 1 N1 7.498u
Rdc1 N1 4 6.2m
Cp1 1 4 7.178p
Rp1 1 4 2854
L2 2 N2 7.498u
Rdc2  N2 3 6.2m
Cp2 2 3 7.178p
Rp2 2 3 2854
Rg1 1 0 500meg
Rg2 2 0 500meg
Rg3 3 0 500meg
Rg4 4 0 500meg
.ends
*******
.subckt 1521_74441521100_10u 1 2 3 4
L1 1 N1 9.098u
Rdc1 N1 4 6.3m
Cp1 1 4 7.474p
Rp1 1 4 2870
L2 2 N2 9.098u
Rdc2  N2 3 6.3m
Cp2 2 3 7.474p
Rp2 2 3 2870
Rg1 1 0 500meg
Rg2 2 0 500meg
Rg3 3 0 500meg
Rg4 4 0 500meg
.ends
*******
.subckt 1521_74441521150_15u 1 2 3 4
L1 1 N1 14.504u
Rdc1 N1 4 8.5m
Cp1 1 4 7.06p
Rp1 1 4 3720
L2 2 N2 14.504u
Rdc2  N2 3 8.5m
Cp2 2 3 7.06p
Rp2 2 3 3720
Rg1 1 0 500meg
Rg2 2 0 500meg
Rg3 3 0 500meg
Rg4 4 0 500meg
.ends
*******
.subckt 1521_74441521220_22u 1 2 3 4
L1 1 N1 21.78u
Rdc1 N1 4 13.6m
Cp1 1 4 7.729p
Rp1 1 4 5558
L2 2 N2 21.78u
Rdc2  N2 3 13.6m
Cp2 2 3 7.729p
Rp2 2 3 5558
Rg1 1 0 500meg
Rg2 2 0 500meg
Rg3 3 0 500meg
Rg4 4 0 500meg
.ends

