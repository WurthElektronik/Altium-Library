**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Aluminum Electrolytic Capacitors
* Matchcode:              WCAP-AI3H
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-30
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 861140783006_2.2mF 1 2
Rser 1 3 0.0256230550864
Lser 2 4 2.7194189038E-08
C1 3 4 0.0022
Rpar 3 4 56407.6392059953
.ends 861140783006_2.2mF
*****
.subckt 861140784012_3.3mF 1 2
Rser 1 3 0.0218909214992
Lser 2 4 3.4460218311E-08
C1 3 4 0.0033
Rpar 3 4 46056.671637863
.ends 861140784012_3.3mF
*****
.subckt 861140786018_4.7mF 1 2
Rser 1 3 0.0240773817871
Lser 2 4 2.0412184406E-08
C1 3 4 0.0047
Rpar 3 4 38592.2999173022
.ends 861140786018_4.7mF
*****
.subckt 861141084008_0.47mF 1 2
Rser 1 3 0.135221660912
Lser 2 4 2.1539930535E-08
C1 3 4 0.00047
Rpar 3 4 217443.301659092
.ends 861141084008_0.47mF
*****
.subckt 861141085015_0.68mF 1 2
Rser 1 3 0.0927957627927
Lser 2 4 2.5557844115E-08
C1 3 4 0.00068
Rpar 3 4 180774.619243458
.ends 861141085015_0.68mF
*****
.subckt 861141085021_1mF 1 2
Rser 1 3 0.0611790824989
Lser 2 4 1.9554137513E-08
C1 3 4 0.001
Rpar 3 4 149071.285888912
.ends 861141085021_1mF
*****
.subckt 861141386015_0.22mF 1 2
Rser 1 3 0.24492
Lser 2 4 1.2918198881E-08
C1 3 4 0.00022
Rpar 3 4 449468.503494618
.ends 861141386015_0.22mF
*****
.subckt 861141386025_0.47mF 1 2
Rser 1 3 0.13499
Lser 2 4 1.3582138314E-08
C1 3 4 0.00047
Rpar 3 4 307510.167054898
.ends 861141386025_0.47mF
*****
.subckt 861141386028_1mF 1 2
Rser 1 3 0.128998276853
Lser 2 4 2.1197282742E-08
C1 3 4 0.001
Rpar 3 4 210818.132467574
.ends 861141386028_1mF
*****
.subckt 861141483001_68uF 1 2
Rser 1 3 0.344
Lser 2 4 1.4759407699E-08
C1 3 4 0.000068
Rpar 3 4 857485.851483451
.ends 861141483001_68uF
*****
.subckt 861141483002_82uF 1 2
Rser 1 3 0.306
Lser 2 4 1.3728290245E-08
C1 3 4 0.000082
Rpar 3 4 780870.410217256
.ends 861141483002_82uF
*****
.subckt 861141483003_0.1mF 1 2
Rser 1 3 0.242
Lser 2 4 1.3346323523E-08
C1 3 4 0.0001
Rpar 3 4 707102.451288498
.ends 861141483003_0.1mF
*****
.subckt 861141483004_0.12mF 1 2
Rser 1 3 0.238
Lser 2 4 1.2778717242E-08
C1 3 4 0.00012
Rpar 3 4 645494.448747741
.ends 861141483004_0.12mF
*****
.subckt 861141483005_0.15mF 1 2
Rser 1 3 0.182
Lser 2 4 1.2725375613E-08
C1 3 4 0.00015
Rpar 3 4 577352.390238896
.ends 861141483005_0.15mF
*****
.subckt 861141483006_0.18mF 1 2
Rser 1 3 0.158
Lser 2 4 1.2711408298E-08
C1 3 4 0.00018
Rpar 3 4 527049.343530762
.ends 861141483006_0.18mF
*****
.subckt 861141483007_0.22mF 1 2
Rser 1 3 0.139
Lser 2 4 1.295154206E-08
C1 3 4 0.00022
Rpar 3 4 476730.266015488
.ends 861141483007_0.22mF
*****
.subckt 861141484008_82uF 1 2
Rser 1 3 0.303
Lser 2 4 1.4951795627E-08
C1 3 4 0.000082
Rpar 3 4 780870.410217256
.ends 861141484008_82uF
*****
.subckt 861141484009_0.1mF 1 2
Rser 1 3 0.274
Lser 2 4 1.4932425828E-08
C1 3 4 0.0001
Rpar 3 4 707102.451288498
.ends 861141484009_0.1mF
*****
.subckt 861141484010_0.12mF 1 2
Rser 1 3 0.244
Lser 2 4 1.4639549587E-08
C1 3 4 0.00012
Rpar 3 4 645494.448747741
.ends 861141484010_0.12mF
*****
.subckt 861141484011_0.15mF 1 2
Rser 1 3 0.195
Lser 2 4 1.3995867639E-08
C1 3 4 0.00015
Rpar 3 4 577352.390238896
.ends 861141484011_0.15mF
*****
.subckt 861141484012_0.18mF 1 2
Rser 1 3 0.178
Lser 2 4 1.3987619065E-08
C1 3 4 0.00018
Rpar 3 4 527049.343530762
.ends 861141484012_0.18mF
*****
.subckt 861141484013_0.22mF 1 2
Rser 1 3 0.12
Lser 2 4 7.78902235300046E-09
C1 3 4 0.00022
Rpar 3 4 476730.266015488
.ends 861141484013_0.22mF
*****
.subckt 861141485014_0.12mF 1 2
Rser 1 3 0.24
Lser 2 4 1.6161837516E-08
C1 3 4 0.00012
Rpar 3 4 645494.448747741
.ends 861141485014_0.12mF
*****
.subckt 861141485015_0.15mF 1 2
Rser 1 3 0.197
Lser 2 4 2.38128565238662E-08
C1 3 4 0.00015
Rpar 3 4 577352.390238896
.ends 861141485015_0.15mF
*****
.subckt 861141485016_0.18mF 1 2
Rser 1 3 0.205
Lser 2 4 2.22199104543036E-08
C1 3 4 0.00018
Rpar 3 4 527049.343530762
.ends 861141485016_0.18mF
*****
.subckt 861141485017_0.22mF 1 2
Rser 1 3 0.154
Lser 2 4 8.82171732329988E-09
C1 3 4 0.00022
Rpar 3 4 476730.266015488
.ends 861141485017_0.22mF
*****
.subckt 861141485018_0.27mF 1 2
Rser 1 3 0.126
Lser 2 4 1.10487045727914E-08
C1 3 4 0.00027
Rpar 3 4 430329.632498494
.ends 861141485018_0.27mF
*****
.subckt 861141485019_0.33mF 1 2
Rser 1 3 0.11
Lser 2 4 9.42208107791878E-09
C1 3 4 0.00033
Rpar 3 4 389249.785912618
.ends 861141485019_0.33mF
*****
.subckt 861141486020_0.22mF 1 2
Rser 1 3 0.142
Lser 2 4 1.3959636387E-08
C1 3 4 0.00022
Rpar 3 4 476730.266015488
.ends 861141486020_0.22mF
*****
.subckt 861141486021_0.27mF 1 2
Rser 1 3 0.117
Lser 2 4 7.96265958601893E-09
C1 3 4 0.00027
Rpar 3 4 430329.632498494
.ends 861141486021_0.27mF
*****
.subckt 861141486022_0.33mF 1 2
Rser 1 3 0.104
Lser 2 4 2.42311788621081E-08
C1 3 4 0.00033
Rpar 3 4 389249.785912618
.ends 861141486022_0.33mF
*****
.subckt 861141486023_0.39mF 1 2
Rser 1 3 0.094
Lser 2 4 2.47745591408481E-08
C1 3 4 0.00039
Rpar 3 4 358057.893983036
.ends 861141486023_0.39mF
*****
.subckt 861141486024_0.47mF 1 2
Rser 1 3 0.085
Lser 2 4 9.61067287881989E-09
C1 3 4 0.00047
Rpar 3 4 326164.952488639
.ends 861141486024_0.47mF
*****
.subckt 861141486025_0.56mF 1 2
Rser 1 3 0.073
Lser 2 4 1.05197206782987E-08
C1 3 4 0.00056
Rpar 3 4 298806.764985159
.ends 861141486025_0.56mF
*****
.subckt 861141486026_0.68mF 1 2
Rser 1 3 0.06
Lser 2 4 1.05528512515298E-08
C1 3 4 0.00068
Rpar 3 4 271162.745854223
.ends 861141486026_0.68mF
*****
.subckt 861140786024_10mF 1 2
Rser 1 3 0.01748
Lser 2 4 1.5255E-08
C1 3 4 10m
Rpar 3 4 124.444
.ends 861140786024_10mF
*****
.subckt 861141485033_470uF  1  2
Rser  1  3   0.086
Lser  2  4  0.000000008
C  3  4  0.00047
Rpar  3  4  326000
.ends  861141485033_470uF
******

















