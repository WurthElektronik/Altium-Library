**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  SMT EMI Suppression Ferrite Bead
* Matchcode:              WE-CBF
* Library Type:           LTspice
* Version:                rev21a
* Created/modified by:    Ella
* Date and Time:          6/18/2024
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2024 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 0402_74279270_40ohm 1 2
Rp 1 2 60
Cp 1 2 0.36p
Rs 1 N3 0.3
L1 N3 2 0.151u
.ends 0402_74279270_40ohm
*******
.subckt 0402_742792701_10ohm 1 2
Rp 1 2 11
Cp 1 2 3.2p
Rs 1 N3 0.05
L1 N3 2 0.04u
.ends 0402_742792701_10ohm
*******
.subckt 0402_74279271_120ohm 1 2
Rp 1 2 182
Cp 1 2 0.343p
Rs 1 N3 0.2
L1 N3 2 0.505u
.ends 0402_74279271_120ohm
*******
.subckt 0402_742792711_100ohm 1 2
Rp 1 2 159
Cp 1 2 0.38p
Rs 1 N3 0.3
L1 N3 2 0.22u
.ends 0402_742792711_100ohm
*******
.subckt 0402_7427927110_10ohm 1 2
Rp 1 2 13
Cp 1 2 1.6p
Rs 1 N3 0.05
L1 N3 2 0.022u
.ends 0402_7427927110_10ohm
*******
.subckt 0402_7427927112_120ohm 1 2
Rp 1 2 850
Cp 1 2 0.337p
Rs 1 N3 0.35
L1 N3 2 0.2u
.ends 0402_7427927112_120ohm
*******
.subckt 0402_7427927115_150ohm 1 2
Rp 1 2 163
Cp 1 2 0.36p
Rs 1 N3 0.4
L1 N3 2 0.27u
.ends 0402_7427927115_150ohm
*******
.subckt 0402_7427927121_220ohm 1 2
Rp 1 2 1510
Cp 1 2 0.405p
Rs 1 N3 0.8
L1 N3 2 0.36u
.ends 0402_7427927121_220ohm
*******
.subckt 0402_7427927130_30ohm 1 2
Rp 1 2 13
Cp 1 2 2.4p
Rs 1 N3 0.15
L1 N3 2 0.025u
.ends 0402_7427927130_30ohm
*******
.subckt 0402_7427927140_47ohm 1 2
Rp 1 2 65
Cp 1 2 0.54p
Rs 1 N3 0.4
L1 N3 2 0.092u
.ends 0402_7427927140_47ohm
*******
.subckt 0402_7427927141_470ohm 1 2
Rp 1 2 1240
Cp 1 2 0.374p
Rs 1 N3 0.45
L1 N3 2 0.73u
.ends 0402_7427927141_470ohm
*******
.subckt 0402_742792716_60ohm 1 2
Rp 1 2 145
Cp 1 2 0.33p
Rs 1 N3 0.25
L1 N3 2 0.985u
.ends 0402_742792716_60ohm
*******
.subckt 0402_7427927160_60ohm 1 2
Rp 1 2 930
Cp 1 2 0.54p
Rs 1 N3 0.3
L1 N3 2 1.6u
.ends 0402_7427927160_60ohm
*******
.subckt 0402_7427927161_600ohm 1 2
Rp 1 2 1300
Cp 1 2 0.38p
Rs 1 N3 0.56
L1 N3 2 0.77u
.ends 0402_7427927161_600ohm
*******
.subckt 0402_7427927170_75ohm 1 2
Rp 1 2 655
Cp 1 2 0.6p
Rs 1 N3 0.31
L1 N3 2 0.12u
.ends 0402_7427927170_75ohm
*******
.subckt 0402_74279272_300ohm 1 2
Rp 1 2 332
Cp 1 2 0.316p
Rs 1 N3 0.8
L1 N3 2 0.076u
.ends 0402_74279272_300ohm
*******
.subckt 0402_7427927218_180ohm 1 2
Rp 1 2 230
Cp 1 2 0.288p
Rs 1 N3 0.3
L1 N3 2 0.39u
.ends 0402_7427927218_180ohm
*******
.subckt 0402_7427927241_470ohm 1 2
Rp 1 2 620
Cp 1 2 0.35p
Rs 1 N3 0.65
L1 N3 2 2u
.ends 0402_7427927241_470ohm
*******
.subckt 0402_7427927261_600ohm 1 2
Rp 1 2 760
Cp 1 2 0.56p
Rs 1 N3 0.6
L1 N3 2 1.15u
.ends 0402_7427927261_600ohm
*******
.subckt 0402_7427927280_80ohm 1 2
Rp 1 2 135
Cp 1 2 0.4p
Rs 1 N3 0.25
L1 N3 2 0.17u
.ends 0402_7427927280_80ohm
*******
.subckt 0402_7427927281_800ohm 1 2
Rp 1 2 530
Cp 1 2 0.36p
Rs 1 N3 0.8
L1 N3 2 1.4u
.ends 0402_7427927281_800ohm
*******
.subckt 0402_7427927291_600ohm 1 2
Rp 1 2 570
Cp 1 2 0.36p
Rs 1 N3 0.6
L1 N3 2 1.6u
.ends 0402_7427927291_600ohm
*******
.subckt 0402_74279273_20ohm 1 2
Rp 1 2 24
Cp 1 2 0.348p
Rs 1 N3 0.2
L1 N3 2 0.622u
.ends 0402_74279273_20ohm
*******
.subckt 0402_742792731_100ohm 1 2
Rp 1 2 130
Cp 1 2 0.38p
Rs 1 N3 0.09
L1 N3 2 0.26u
.ends 0402_742792731_100ohm
*******
.subckt 0402_7427927310_10ohm 1 2
Rp 1 2 12
Cp 1 2 2p
Rs 1 N3 0.03
L1 N3 2 0.033u
.ends 0402_7427927310_10ohm
*******
.subckt 0402_7427927311_120ohm 1 2
Rp 1 2 135
Cp 1 2 0.3p
Rs 1 N3 0.09
L1 N3 2 0.3u
.ends 0402_7427927311_120ohm
*******
.subckt 0402_7427927370_70ohm 1 2
Rp 1 2 73
Cp 1 2 0.38p
Rs 1 N3 0.09
L1 N3 2 0.178u
.ends 0402_7427927370_70ohm
*******
.subckt 0402_74279274_30ohm 1 2
Rp 1 2 39
Cp 1 2 0.266p
Rs 1 N3 0.25
L1 N3 2 0.108u
.ends 0402_74279274_30ohm
*******
.subckt 0402_74279276_60ohm 1 2
Rp 1 2 103
Cp 1 2 0.273p
Rs 1 N3 0.35
L1 N3 2 0.192u
.ends 0402_74279276_60ohm
*******
.subckt 0402_74279277_70ohm 1 2
Rp 1 2 102
Cp 1 2 0.255p
Rs 1 N3 0.15
L1 N3 2 0.273u
.ends 0402_74279277_70ohm
*******
.subckt 0402_74279278_240ohm 1 2
Rp 1 2 361
Cp 1 2 0.275p
Rs 1 N3 0.7
L1 N3 2 0.911u
.ends 0402_74279278_240ohm
*******
.subckt 0402_742792780_220ohm 1 2
Rp 1 2 270
Cp 1 2 0.42p
Rs 1 N3 0.35
L1 N3 2 0.67u
.ends 0402_742792780_220ohm
*******
.subckt 0402_74279279_600ohm 1 2
Rp 1 2 785
Cp 1 2 0.535p
Rs 1 N3 1
L1 N3 2 1.545u
.ends 0402_74279279_600ohm
*******
.subckt 0402_742792796_1000ohm 1 2
Rp 1 2 1100
Cp 1 2 0.58p
Rs 1 N3 1.5
L1 N3 2 2.6u
.ends 0402_742792796_1000ohm
*******
.subckt 0603_74279260_40ohm 1 2
Rp 1 2 85
Cp 1 2 0.212p
Rs 1 N3 0.15
L1 N3 2 0.104u
.ends 0603_74279260_40ohm
*******
.subckt 0603_742792601_30ohm 1 2
Rp 1 2 51
Cp 1 2 0.092p
Rs 1 N3 0.03
L1 N3 2 0.073u
.ends 0603_742792601_30ohm
*******
.subckt 0603_742792602_60ohm 1 2
Rp 1 2 90
Cp 1 2 0.275p
Rs 1 N3 0.04
L1 N3 2 0.148u
.ends 0603_742792602_60ohm
*******
.subckt 0603_742792603_28ohm 1 2
Rp 1 2 44
Cp 1 2 0.144p
Rs 1 N3 0.03
L1 N3 2 0.068u
.ends 0603_742792603_28ohm
*******
.subckt 0603_742792604_22ohm 1 2
Rp 1 2 42
Cp 1 2 0.07p
Rs 1 N3 0.05
L1 N3 2 0.066u
.ends 0603_742792604_22ohm
*******
.subckt 0603_742792605_33ohm 1 2
Rp 1 2 45
Cp 1 2 0.073p
Rs 1 N3 0.1
L1 N3 2 0.07u
.ends 0603_742792605_33ohm
*******
.subckt 0603_742792606_120ohm 1 2
Rp 1 2 500
Cp 1 2 0.8p
Rs 1 N3 0.35
L1 N3 2 0.19u
.ends 0603_742792606_120ohm
*******
.subckt 0603_742792607_68ohm 1 2
Rp 1 2 300
Cp 1 2 0.738p
Rs 1 N3 0.3
L1 N3 2 0.1u
.ends 0603_742792607_68ohm
*******
.subckt 0603_742792608_47ohm 1 2
Rp 1 2 75
Cp 1 2 0.04p
Rs 1 N3 0.1
L1 N3 2 0.1u
.ends 0603_742792608_47ohm
*******
.subckt 0603_742792609_30ohm 1 2
Rp 1 2 35
Cp 1 2 0.85p
Rs 1 N3 0.04
L1 N3 2 0.15u
.ends 0603_742792609_30ohm
*******
.subckt 0603_74279261_80ohm 1 2
Rp 1 2 321
Cp 1 2 0.496p
Rs 1 N3 0.3
L1 N3 2 0.132u
.ends 0603_74279261_80ohm
*******
.subckt 0603_74279262_120ohm 1 2
Rp 1 2 172
Cp 1 2 0.545p
Rs 1 N3 0.3
L1 N3 2 0.37u
.ends 0603_74279262_120ohm
*******
.subckt 0603_742792620_100ohm 1 2
Rp 1 2 120
Cp 1 2 0.68p
Rs 1 N3 0.15
L1 N3 2 0.034u
.ends 0603_742792620_100ohm
*******
.subckt 0603_742792621_140ohm 1 2
Rp 1 2 408
Cp 1 2 0.585p
Rs 1 N3 0.2
L1 N3 2 0.2u
.ends 0603_742792621_140ohm
*******
.subckt 0603_742792622_180ohm 1 2
Rp 1 2 277
Cp 1 2 0.68p
Rs 1 N3 0.3
L1 N3 2 0.434u
.ends 0603_742792622_180ohm
*******
.subckt 0603_742792624_180ohm 1 2
Rp 1 2 260
Cp 1 2 0.67p
Rs 1 N3 0.09
L1 N3 2 0.42u
.ends 0603_742792624_180ohm
*******
.subckt 0603_742792625_120ohm 1 2
Rp 1 2 140
Cp 1 2 0.56p
Rs 1 N3 0.05
L1 N3 2 0.325u
.ends 0603_742792625_120ohm
*******
.subckt 0603_74279263_220ohm 1 2
Rp 1 2 330
Cp 1 2 0.49p
Rs 1 N3 0.3
L1 N3 2 0.523u
.ends 0603_74279263_220ohm
*******
.subckt 0603_742792631_240ohm 1 2
Rp 1 2 384
Cp 1 2 0.56p
Rs 1 N3 0.4
L1 N3 2 0.67u
.ends 0603_742792631_240ohm
*******
.subckt 0603_74279264_300ohm 1 2
Rp 1 2 484
Cp 1 2 0.48p
Rs 1 N3 0.35
L1 N3 2 0.516u
.ends 0603_74279264_300ohm
*******
.subckt 0603_742792640_300ohm 1 2
Rp 1 2 1950
Cp 1 2 0.8p
Rs 1 N3 0.35
L1 N3 2 0.47u
.ends 0603_742792640_300ohm
*******
.subckt 0603_742792641_300ohm 1 2
Rp 1 2 503
Cp 1 2 0.462p
Rs 1 N3 0.15
L1 N3 2 0.782u
.ends 0603_742792641_300ohm
*******
.subckt 0603_742792642_470ohm 1 2
Rp 1 2 662
Cp 1 2 0.608p
Rs 1 N3 0.45
L1 N3 2 1.164u
.ends 0603_742792642_470ohm
*******
.subckt 0603_742792643_470ohm 1 2
Rp 1 2 810
Cp 1 2 0.76p
Rs 1 N3 0.35
L1 N3 2 0.7u
.ends 0603_742792643_470ohm
*******
.subckt 0603_742792645_470ohm 1 2
Rp 1 2 420
Cp 1 2 0.7p
Rs 1 N3 0.2
L1 N3 2 1.3u
.ends 0603_742792645_470ohm
*******
.subckt 0603_74279265_600ohm 1 2
Rp 1 2 752
Cp 1 2 0.67p
Rs 1 N3 0.45
L1 N3 2 1.8u
.ends 0603_74279265_600ohm
*******
.subckt 0603_742792651_600ohm 1 2
Rp 1 2 813
Cp 1 2 0.617p
Rs 1 N3 0.2
L1 N3 2 1.384u
.ends 0603_742792651_600ohm
*******
.subckt 0603_742792653_600ohm 1 2
Rp 1 2 5400
Cp 1 2 1p
Rs 1 N3 0.65
L1 N3 2 0.68u
.ends 0603_742792653_600ohm
*******
.subckt 0603_742792656_750ohm 1 2
Rp 1 2 790
Cp 1 2 0.78p
Rs 1 N3 0.35
L1 N3 2 2.6u
.ends 0603_742792656_750ohm
*******
.subckt 0603_74279266_1000ohm 1 2
Rp 1 2 1290
Cp 1 2 0.604p
Rs 1 N3 0.6
L1 N3 2 2.393u
.ends 0603_74279266_1000ohm
*******
.subckt 0603_742792662_1000ohm 1 2
Rp 1 2 1050
Cp 1 2 0.68p
Rs 1 N3 0.3
L1 N3 2 3.3u
.ends 0603_742792662_1000ohm
*******
.subckt 0603_742792663_1000ohm 1 2
Rp 1 2 1320
Cp 1 2 0.57p
Rs 1 N3 0.85
L1 N3 2 1.45u
.ends 0603_742792663_1000ohm
*******
.subckt 0603_742792664_1000ohm 1 2
Rp 1 2 1800
Cp 1 2 0.79p
Rs 1 N3 0.6
L1 N3 2 1.16u
.ends 0603_742792664_1000ohm
*******
.subckt 0603_74279267_60ohm 1 2
Rp 1 2 75
Cp 1 2 0.25p
Rs 1 N3 0.3
L1 N3 2 0.258u
.ends 0603_74279267_60ohm
*******
.subckt 0603_74279268_15ohm 1 2
Rp 1 2 78
Cp 1 2 0.256p
Rs 1 N3 0.1
L1 N3 2 0.021u
.ends 0603_74279268_15ohm
*******
.subckt 0603_74279269_1200ohm 1 2
Rp 1 2 1336
Cp 1 2 0.622p
Rs 1 N3 0.7
L1 N3 2 2.583u
.ends 0603_74279269_1200ohm
*******
.subckt 0603_742792691_1500ohm 1 2
Rp 1 2 1817
Cp 1 2 0.808p
Rs 1 N3 0.7
L1 N3 2 3.08u
.ends 0603_742792691_1500ohm
*******
.subckt 0603_742792692_1800ohm 1 2
Rp 1 2 1940
Cp 1 2 0.672p
Rs 1 N3 0.8
L1 N3 2 2.4u
.ends 0603_742792692_1800ohm
*******
.subckt 0603_742792693_2200ohm 1 2
Rp 1 2 2054
Cp 1 2 0.911p
Rs 1 N3 0.8
L1 N3 2 2.58u
.ends 0603_742792693_2200ohm
*******
.subckt 0603_742792695_2500ohm 1 2
Rp 1 2 2600
Cp 1 2 0.73p
Rs 1 N3 1
L1 N3 2 2.7u
.ends 0603_742792695_2500ohm
*******
.subckt 0805_7427920_11ohm 1 2
Rp 1 2 19
Cp 1 2 0.235p
Rs 1 N3 0.15
L1 N3 2 0.016u
.ends 0805_7427920_11ohm
*******
.subckt 0805_742792005_5ohm 1 2
Rp 1 2 14
Cp 1 2 0.5p
Rs 1 N3 0.07
L1 N3 2 0.075u
.ends 0805_742792005_5ohm
*******
.subckt 0805_74279201_32ohm 1 2
Rp 1 2 70
Cp 1 2 0.178p
Rs 1 N3 0.15
L1 N3 2 0.054u
.ends 0805_74279201_32ohm
*******
.subckt 0805_742792010_7ohm 1 2
Rp 1 2 12
Cp 1 2 0.001p
Rs 1 N3 0.03
L1 N3 2 0.018u
.ends 0805_742792010_7ohm
*******
.subckt 0805_742792011_10ohm 1 2
Rp 1 2 23
Cp 1 2 0.241p
Rs 1 N3 0.025
L1 N3 2 0.023u
.ends 0805_742792011_10ohm
*******
.subckt 0805_742792012_33ohm 1 2
Rp 1 2 80
Cp 1 2 0.067p
Rs 1 N3 0.008
L1 N3 2 0.093u
.ends 0805_742792012_33ohm
*******
.subckt 0805_742792015_56ohm 1 2
Rp 1 2 260
Cp 1 2 0.667p
Rs 1 N3 0.3
L1 N3 2 0.089u
.ends 0805_742792015_56ohm
*******
.subckt 0805_742792017_90ohm 1 2
Rp 1 2 135
Cp 1 2 0.465p
Rs 1 N3 0.02
L1 N3 2 0.26u
.ends 0805_742792017_90ohm
*******
.subckt 0805_74279202_120ohm 1 2
Rp 1 2 170
Cp 1 2 0.831p
Rs 1 N3 0.1
L1 N3 2 0.35u
.ends 0805_74279202_120ohm
*******
.subckt 0805_742792021_22ohm 1 2
Rp 1 2 37
Cp 1 2 0.275p
Rs 1 N3 0.008
L1 N3 2 0.047u
.ends 0805_742792021_22ohm
*******
.subckt 0805_742792022_220ohm 1 2
Rp 1 2 360
Cp 1 2 0.68p
Rs 1 N3 0.05
L1 N3 2 0.564u
.ends 0805_742792022_220ohm
*******
.subckt 0805_742792023_120ohm 1 2
Rp 1 2 177
Cp 1 2 0.847p
Rs 1 N3 0.03
L1 N3 2 0.377u
.ends 0805_742792023_120ohm
*******
.subckt 0805_742792025_120ohm 1 2
Rp 1 2 145
Cp 1 2 0.95p
Rs 1 N3 0.02
L1 N3 2 0.197u
.ends 0805_742792025_120ohm
*******
.subckt 0805_74279203_150ohm 1 2
Rp 1 2 240
Cp 1 2 0.812p
Rs 1 N3 0.25
L1 N3 2 0.364u
.ends 0805_74279203_150ohm
*******
.subckt 0805_742792030_30ohm 1 2
Rp 1 2 39
Cp 1 2 0.75p
Rs 1 N3 0.003
L1 N3 2 0.059u
.ends 0805_742792030_30ohm
*******
.subckt 0805_742792031_300ohm 1 2
Rp 1 2 330
Cp 1 2 1.12p
Rs 1 N3 0.05
L1 N3 2 1.21u
.ends 0805_742792031_300ohm
*******
.subckt 0805_742792032_400ohm 1 2
Rp 1 2 495
Cp 1 2 1.25p
Rs 1 N3 0.3
L1 N3 2 2.07u
.ends 0805_742792032_400ohm
*******
.subckt 0805_742792034_220ohm 1 2
Rp 1 2 352
Cp 1 2 0.664p
Rs 1 N3 0.3
L1 N3 2 0.563u
.ends 0805_742792034_220ohm
*******
.subckt 0805_742792035_300ohm 1 2
Rp 1 2 430
Cp 1 2 0.855p
Rs 1 N3 0.3
L1 N3 2 0.448u
.ends 0805_742792035_300ohm
*******
.subckt 0805_742792036_470ohm 1 2
Rp 1 2 559
Cp 1 2 0.884p
Rs 1 N3 0.3
L1 N3 2 1.018u
.ends 0805_742792036_470ohm
*******
.subckt 0805_742792037_330ohm 1 2
Rp 1 2 362
Cp 1 2 0.863p
Rs 1 N3 0.08
L1 N3 2 0.775u
.ends 0805_742792037_330ohm
*******
.subckt 0805_742792038_240ohm 1 2
Rp 1 2 302
Cp 1 2 1.5p
Rs 1 N3 0.4
L1 N3 2 0.435u
.ends 0805_742792038_240ohm
*******
.subckt 0805_74279204_600ohm 1 2
Rp 1 2 754
Cp 1 2 0.784p
Rs 1 N3 0.35
L1 N3 2 1.381u
.ends 0805_74279204_600ohm
*******
.subckt 0805_742792040_600ohm 1 2
Rp 1 2 830
Cp 1 2 0.836p
Rs 1 N3 0.15
L1 N3 2 1.43u
.ends 0805_742792040_600ohm
*******
.subckt 0805_742792041_600ohm 1 2
Rp 1 2 730
Cp 1 2 0.791p
Rs 1 N3 0.4
L1 N3 2 1.2u
.ends 0805_742792041_600ohm
*******
.subckt 0805_7427920415_600ohm 1 2
Rp 1 2 540
Cp 1 2 1.04p
Rs 1 N3 0.3
L1 N3 2 2.6u
.ends 0805_7427920415_600ohm
*******
.subckt 0805_742792042_600ohm 1 2
Rp 1 2 3380
Cp 1 2 1.1p
Rs 1 N3 0.5
L1 N3 2 0.7u
.ends 0805_742792042_600ohm
*******
.subckt 0805_742792043_600ohm 1 2
Rp 1 2 6300
Cp 1 2 1.2p
Rs 1 N3 0.65
L1 N3 2 0.61u
.ends 0805_742792043_600ohm
*******
.subckt 0805_742792045_750ohm 1 2
Rp 1 2 1080
Cp 1 2 1.1p
Rs 1 N3 0.3
L1 N3 2 0.89u
.ends 0805_742792045_750ohm
*******
.subckt 0805_74279205_1000ohm 1 2
Rp 1 2 1198
Cp 1 2 0.853p
Rs 1 N3 0.45
L1 N3 2 2u
.ends 0805_74279205_1000ohm
*******
.subckt 0805_74279206_30ohm 1 2
Rp 1 2 59
Cp 1 2 0.2p
Rs 1 N3 0.025
L1 N3 2 0.08u
.ends 0805_74279206_30ohm
*******
.subckt 0805_742792062_80ohm 1 2
Rp 1 2 137
Cp 1 2 0.306p
Rs 1 N3 0.2
L1 N3 2 0.138u
.ends 0805_742792062_80ohm
*******
.subckt 0805_742792063_60ohm 1 2
Rp 1 2 100
Cp 1 2 0.712p
Rs 1 N3 0.025
L1 N3 2 0.141u
.ends 0805_742792063_60ohm
*******
.subckt 0805_742792064_75ohm 1 2
Rp 1 2 270
Cp 1 2 0.931p
Rs 1 N3 0.2
L1 N3 2 0.128u
.ends 0805_742792064_75ohm
*******
.subckt 0805_74279207_100ohm 1 2
Rp 1 2 220
Cp 1 2 0.526p
Rs 1 N3 0.15
L1 N3 2 0.25u
.ends 0805_74279207_100ohm
*******
.subckt 0805_74279208_40ohm 1 2
Rp 1 2 64
Cp 1 2 0.1p
Rs 1 N3 0.15
L1 N3 2 0.08u
.ends 0805_74279208_40ohm
*******
.subckt 0805_74279209_1200ohm 1 2
Rp 1 2 1458
Cp 1 2 0.986p
Rs 1 N3 0.55
L1 N3 2 1.47u
.ends 0805_74279209_1200ohm
*******
.subckt 0805_742792090_1800ohm 1 2
Rp 1 2 2350
Cp 1 2 1.2p
Rs 1 N3 0.4
L1 N3 2 1.4u
.ends 0805_742792090_1800ohm
*******
.subckt 0805_742792091_1500ohm 1 2
Rp 1 2 1500
Cp 1 2 1.04p
Rs 1 N3 0.55
L1 N3 2 1.385u
.ends 0805_742792091_1500ohm
*******
.subckt 0805_742792092_2000ohm 1 2
Rp 1 2 2700
Cp 1 2 1.122p
Rs 1 N3 0.6
L1 N3 2 3.642u
.ends 0805_742792092_2000ohm
*******
.subckt 0805_742792093_2200ohm 1 2
Rp 1 2 2780
Cp 1 2 0.97p
Rs 1 N3 0.6
L1 N3 2 3.42u
.ends 0805_742792093_2200ohm
*******
.subckt 0805_742792094_2200ohm 1 2
Rp 1 2 2500
Cp 1 2 1.2p
Rs 1 N3 0.5
L1 N3 2 1.3u
.ends 0805_742792094_2200ohm
*******
.subckt 0805_742792095_2700ohm 1 2
Rp 1 2 3700
Cp 1 2 1.4p
Rs 1 N3 0.6
L1 N3 2 1.5u
.ends 0805_742792095_2700ohm
*******
.subckt 0805_742792096_1000ohm 1 2
Rp 1 2 1080
Cp 1 2 1.3p
Rs 1 N3 0.3
L1 N3 2 5.3u
.ends 0805_742792096_1000ohm
*******
.subckt 0805_742792097_1500ohm 1 2
Rp 1 2 1570
Cp 1 2 1.34p
Rs 1 N3 0.3
L1 N3 2 8.3u
.ends 0805_742792097_1500ohm
*******
.subckt 1206_7427921_32ohm 1 2
Rp 1 2 53
Cp 1 2 0.235p
Rs 1 N3 0.2
L1 N3 2 0.086u
.ends 1206_7427921_32ohm
*******
.subckt 1206_74279210_30ohm 1 2
Rp 1 2 51
Cp 1 2 0.024p
Rs 1 N3 0.04
L1 N3 2 0.075u
.ends 1206_74279210_30ohm
*******
.subckt 1206_74279211_90ohm 1 2
Rp 1 2 256
Cp 1 2 0.274p
Rs 1 N3 0.3
L1 N3 2 0.204u
.ends 1206_74279211_90ohm
*******
.subckt 1206_742792110_19ohm 1 2
Rp 1 2 90
Cp 1 2 0.001p
Rs 1 N3 0.04
L1 N3 2 0.029u
.ends 1206_742792110_19ohm
*******
.subckt 1206_742792111_26ohm 1 2
Rp 1 2 30
Cp 1 2 0.001p
Rs 1 N3 0.04
L1 N3 2 0.09u
.ends 1206_742792111_26ohm
*******
.subckt 1206_742792112_31ohm 1 2
Rp 1 2 56
Cp 1 2 0.197p
Rs 1 N3 0.04
L1 N3 2 0.064u
.ends 1206_742792112_31ohm
*******
.subckt 1206_742792113_120ohm 1 2
Rp 1 2 160
Cp 1 2 0.605p
Rs 1 N3 0.03
L1 N3 2 0.404u
.ends 1206_742792113_120ohm
*******
.subckt 1206_742792114_50ohm 1 2
Rp 1 2 52
Cp 1 2 0.04p
Rs 1 N3 0.025
L1 N3 2 0.145u
.ends 1206_742792114_50ohm
*******
.subckt 1206_742792115_80ohm 1 2
Rp 1 2 122
Cp 1 2 0.312p
Rs 1 N3 0.025
L1 N3 2 0.2u
.ends 1206_742792115_80ohm
*******
.subckt 1206_742792116_500ohm 1 2
Rp 1 2 550
Cp 1 2 1.179p
Rs 1 N3 0.06
L1 N3 2 1.62u
.ends 1206_742792116_500ohm
*******
.subckt 1206_742792117_48ohm 1 2
Rp 1 2 73
Cp 1 2 0.083p
Rs 1 N3 0.005
L1 N3 2 0.084u
.ends 1206_742792117_48ohm
*******
.subckt 1206_742792118_600ohm 1 2
Rp 1 2 620
Cp 1 2 1.9p
Rs 1 N3 0.07
L1 N3 2 1.8u
.ends 1206_742792118_600ohm
*******
.subckt 1206_742792121_300ohm 1 2
Rp 1 2 290
Cp 1 2 1.45p
Rs 1 N3 0.06
L1 N3 2 0.95u
.ends 1206_742792121_300ohm
*******
.subckt 1206_742792122_220ohm 1 2
Rp 1 2 300
Cp 1 2 1.04p
Rs 1 N3 0.3
L1 N3 2 0.54u
.ends 1206_742792122_220ohm
*******
.subckt 1206_742792124_470ohm 1 2
Rp 1 2 540
Cp 1 2 1.928p
Rs 1 N3 0.3
L1 N3 2 1.113u
.ends 1206_742792124_470ohm
*******
.subckt 1206_74279213_600ohm 1 2
Rp 1 2 632
Cp 1 2 1.845p
Rs 1 N3 0.3
L1 N3 2 1.45u
.ends 1206_74279213_600ohm
*******
.subckt 1206_742792131_600ohm 1 2
Rp 1 2 620
Cp 1 2 1.213p
Rs 1 N3 0.3
L1 N3 2 1.267u
.ends 1206_742792131_600ohm
*******
.subckt 1206_742792133_600ohm 1 2
Rp 1 2 910
Cp 1 2 3.103p
Rs 1 N3 0.3
L1 N3 2 1.644u
.ends 1206_742792133_600ohm
*******
.subckt 1206_74279214_1000ohm 1 2
Rp 1 2 1100
Cp 1 2 1.367p
Rs 1 N3 0.45
L1 N3 2 2.074u
.ends 1206_74279214_1000ohm
*******
.subckt 1206_742792141_1000ohm 1 2
Rp 1 2 1050
Cp 1 2 1.145p
Rs 1 N3 0.3
L1 N3 2 4.6u
.ends 1206_742792141_1000ohm
*******
.subckt 1206_74279215_80ohm 1 2
Rp 1 2 94
Cp 1 2 0.16p
Rs 1 N3 0.03
L1 N3 2 0.241u
.ends 1206_74279215_80ohm
*******
.subckt 1206_742792150_80ohm 1 2
Rp 1 2 88
Cp 1 2 0.072p
Rs 1 N3 0.02
L1 N3 2 0.252u
.ends 1206_742792150_80ohm
*******
.subckt 1206_742792151_70ohm 1 2
Rp 1 2 100
Cp 1 2 0.145p
Rs 1 N3 0.3
L1 N3 2 0.223u
.ends 1206_742792151_70ohm
*******
.subckt 1206_74279216_1200ohm 1 2
Rp 1 2 1450
Cp 1 2 1.45p
Rs 1 N3 0.5
L1 N3 2 1.9u
.ends 1206_74279216_1200ohm
*******
.subckt 1206_742792161_1000ohm 1 2
Rp 1 2 1500
Cp 1 2 1.2p
Rs 1 N3 0.5
L1 N3 2 0.0065u
.ends 1206_742792161_1000ohm
*******
.subckt 1206_74279217_1000ohm 1 2
Rp 1 2 2223
Cp 1 2 1.5p
Rs 1 N3 0.45
L1 N3 2 0.0047u
.ends 1206_74279217_1000ohm
*******
.subckt 1206_74279218_600ohm 1 2
Rp 1 2 587
Cp 1 2 1.216p
Rs 1 N3 0.1
L1 N3 2 1.542u
.ends 1206_74279218_600ohm
*******
.subckt 1206_74279219_700ohm 1 2
Rp 1 2 2150
Cp 1 2 1.5p
Rs 1 N3 0.65
L1 N3 2 7.3u
.ends 1206_74279219_700ohm
*******
.subckt 1206_7427922_60ohm 1 2
Rp 1 2 110
Cp 1 2 0.09p
Rs 1 N3 0.2
L1 N3 2 0.11u
.ends 1206_7427922_60ohm
*******
.subckt 1210_7427923_90ohm 1 2
Rp 1 2 207
Cp 1 2 0.247p
Rs 1 N3 0.3
L1 N3 2 0.145u
.ends 1210_7427923_90ohm
*******
.subckt 1210_74279230_32ohm 1 2
Rp 1 2 62
Cp 1 2 0.25p
Rs 1 N3 0.3
L1 N3 2 0.084u
.ends 1210_74279230_32ohm
*******
.subckt 1210_74279231_60ohm 1 2
Rp 1 2 92
Cp 1 2 0.35p
Rs 1 N3 0.3
L1 N3 2 0.12u
.ends 1210_74279231_60ohm
*******
.subckt 1210_742792310_30ohm 1 2
Rp 1 2 62
Cp 1 2 0.242p
Rs 1 N3 0.05
L1 N3 2 0.1u
.ends 1210_742792310_30ohm
*******
.subckt 1210_742792311_52ohm 1 2
Rp 1 2 96
Cp 1 2 0.026p
Rs 1 N3 0.05
L1 N3 2 0.155u
.ends 1210_742792311_52ohm
*******
.subckt 1210_742792312_65ohm 1 2
Rp 1 2 100
Cp 1 2 0.025p
Rs 1 N3 0.03
L1 N3 2 0.14u
.ends 1210_742792312_65ohm
*******
.subckt 1806_7427924_60ohm 1 2
Rp 1 2 125
Cp 1 2 0.056p
Rs 1 N3 0.3
L1 N3 2 0.148u
.ends 1806_7427924_60ohm
*******
.subckt 1806_74279241_80ohm 1 2
Rp 1 2 120
Cp 1 2 0.102p
Rs 1 N3 0.3
L1 N3 2 0.213u
.ends 1806_74279241_80ohm
*******
.subckt 1806_742792410_60ohm 1 2
Rp 1 2 111
Cp 1 2 0.034p
Rs 1 N3 0.01
L1 N3 2 0.148u
.ends 1806_742792410_60ohm
*******
.subckt 1806_742792411_80ohm 1 2
Rp 1 2 80
Cp 1 2 0.04p
Rs 1 N3 0.04
L1 N3 2 0.3u
.ends 1806_742792411_80ohm
*******
.subckt 1806_74279242_150ohm 1 2
Rp 1 2 221
Cp 1 2 0.62p
Rs 1 N3 0.5
L1 N3 2 0.4u
.ends 1806_74279242_150ohm
*******
.subckt 1806_74279243_75ohm 1 2
Rp 1 2 154
Cp 1 2 0.044p
Rs 1 N3 0.025
L1 N3 2 0.18u
.ends 1806_74279243_75ohm
*******
.subckt 1806_74279244_850ohm 1 2
Rp 1 2 1146
Cp 1 2 2.55p
Rs 1 N3 0.1
L1 N3 2 3.541u
.ends 1806_74279244_850ohm
*******
.subckt 1806_74279245_110ohm 1 2
Rp 1 2 145
Cp 1 2 0.006p
Rs 1 N3 0.035
L1 N3 2 0.23u
.ends 1806_74279245_110ohm
*******
.subckt 1806_74279246_1000ohm 1 2
Rp 1 2 1045
Cp 1 2 1.241p
Rs 1 N3 0.056
L1 N3 2 3.003u
.ends 1806_74279246_1000ohm
*******
.subckt 1812_7427925_120ohm 1 2
Rp 1 2 192
Cp 1 2 0.42p
Rs 1 N3 0.3
L1 N3 2 0.293u
.ends 1812_7427925_120ohm
*******
.subckt 1812_74279250_70ohm 1 2
Rp 1 2 100
Cp 1 2 0.067p
Rs 1 N3 0.3
L1 N3 2 0.285u
.ends 1812_74279250_70ohm
*******
.subckt 1812_742792510_70ohm 1 2
Rp 1 2 100
Cp 1 2 0.101p
Rs 1 N3 0.03
L1 N3 2 0.284u
.ends 1812_742792510_70ohm
*******
.subckt 1812_742792511_120ohm 1 2
Rp 1 2 152
Cp 1 2 0.36p
Rs 1 N3 0.05
L1 N3 2 0.482u
.ends 1812_742792511_120ohm
*******
.subckt 1812_742792514_600ohm 1 2
Rp 1 2 981
Cp 1 2 4.9p
Rs 1 N3 0.04
L1 N3 2 1.116u
.ends 1812_742792514_600ohm
*******
.subckt 1812_742792515_785ohm 1 2
Rp 1 2 1616
Cp 1 2 3.6p
Rs 1 N3 0.05
L1 N3 2 1.4u
.ends 1812_742792515_785ohm
*******
.subckt 1812_74279252_880ohm 1 2
Rp 1 2 1012
Cp 1 2 4p
Rs 1 N3 0.035
L1 N3 2 0.633u
.ends 1812_74279252_880ohm
*******
.subckt 2220_7427928101_100Ohm 1 2
Rp 1 2 156.47251
Cp 1 2 0.21122376p
Rs 1 N3 0.004
L1 N3 2 0.221105441u
.ends 2220_7427928101_100Ohm
*******
.subckt 2220_7427928161_160Ohm 1 2
Rp 1 2 242.300464
Cp 1 2 0.233347318p
Rs 1 N3 0.008
L1 N3 2 0.35733144u
.ends 2220_7427928161_160Ohm
*******
.subckt 2220_7427928251_250Ohm 1 2
Rp 1 2 308.804555
Cp 1 2 1.305564p
Rs 1 N3 0.007
L1 N3 2 0.770870664u
.ends 2220_7427928251_250Ohm
*******
.subckt 2220_7427928551_500Ohm 1 2
Rp 1 2 795.422519
Cp 1 2 0.300104809p
Rs 1 N3 0.0023
L1 N3 2 1.294086u
.ends 2220_7427928551_500Ohm
*******
.subckt 2220_7427928601_600Ohm 1 2
Rp 1 2 646.353978
Cp 1 2 2.270116p
Rs 1 N3 0.01
L1 N3 2 1.008701959u
.ends 2220_7427928601_600Ohm
*******
.subckt 2220_7427928801_800Ohm 1 2
Rp 1 2 806.614005
Cp 1 2 2.45024p
Rs 1 N3 0.006
L1 N3 2 0.975124u
.ends 2220_7427928801_800Ohm
*******
