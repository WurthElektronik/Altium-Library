**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Polymer Capacitors
* Matchcode:             WCAP-PHSE
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 875046219001_330uF 1 2
Rser 1 3 0.00194837289123
Lser 2 4 0.000000001
C1 3 4 0.00033
Rpar 3 4 30303.0303030303
.ends 875046219001_330uF
*******
.subckt 875046219002_470uF 1 2
Rser 1 3 0.0015259349176
Lser 2 4 0.00000000049
C1 3 4 0.00047
Rpar 3 4 21276.5957446809
.ends 875046219002_470uF
*******
.subckt 875046219003_560uF 1 2
Rser 1 3 0.00197709932745
Lser 2 4 0.00000000059
C1 3 4 0.00056
Rpar 3 4 17857.1428571429
.ends 875046219003_560uF
*******
.subckt 875046319001_470uF 1 2
Rser 1 3 0.00194601517173
Lser 2 4 0.00000000062
C1 3 4 0.00047
Rpar 3 4 21276.5957446809
.ends 875046319001_470uF
*******
