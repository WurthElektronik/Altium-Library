**************************************************
* Manufacturer:          Würth Elektronik 
* Kinds:                 Multilayer Ceramic Chip Capacitors
* Matchcode:             WCAP-CSST
* Library Type:          LTspice
* Version:               rev24a
* Created/modified by:   Ella
* Date and Time:         7/11/2024
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2024 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************
.subckt 0603_885382206001_220pF 1 2
Rser 1 3 0.0015
Lser 2 4 0.0000000005
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885382206001_220pF
*******
.subckt 0603_885382206002_10nF 1 2
Rser 1 3 0.19
Lser 2 4 8.43227742E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885382206002_10nF
*******
.subckt 0603_885382206003_22nF 1 2
Rser 1 3 0.09
Lser 2 4 8.02867112E-10
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885382206003_22nF
*******
.subckt 0603_885382206004_100nF 1 2
Rser 1 3 0.105
Lser 2 4 7.84352286E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885382206004_100nF
*******
.subckt 0603_885382206005_1nF 1 2
Rser 1 3 0.1
Lser 2 4 7.70337339E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885382206005_1nF
*******
.subckt 0805_885382207001_1uF 1 2
Rser 1 3 0.0237265668732
Lser 2 4 8.71815019E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885382207001_1uF
*******
.subckt 0805_885382207002_330nF 1 2
Rser 1 3 0.053
Lser 2 4 8.98145352E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885382207002_330nF
*******
.subckt 0805_885382207003_1uF 1 2
Rser 1 3 0.020128437829
Lser 2 4 8.47599532E-10
C1 3 4 9.20438317942E-07
Rpar 3 4 500000000
.ends 0805_885382207003_1uF
*******
.subckt 0805_885382207004_1nF 1 2
Rser 1 3 0.11
Lser 2 4 8.48075201E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885382207004_1nF
*******
.subckt 0805_885382207005_2.2nF 1 2
Rser 1 3 0.11
Lser 2 4 9.60090407E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885382207005_2.2nF
*******
.subckt 0805_885382207006_10nF 1 2
Rser 1 3 0.065
Lser 2 4 1.014725274E-09
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885382207006_10nF
*******
.subckt 0805_885382207007_100nF 1 2
Rser 1 3 0.0397714465846
Lser 2 4 9.11116414E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885382207007_100nF
*******
.subckt 0805_885382207008_220nF 1 2
Rser 1 3 0.0518795851536
Lser 2 4 9.05805992E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885382207008_220nF
*******
.subckt 0805_885382207009_10nF 1 2
Rser 1 3 0.0761569081315
Lser 2 4 9.53244591E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885382207009_10nF
*******
.subckt 0805_885382207010_270pF 1 2
Rser 1 3 0.8
Lser 2 4 0.00000000075
C1 3 4 0.00000000027
Rpar 3 4 10000000000
.ends 0805_885382207010_270pF
*******
.subckt 0805_885382207011_1nF 1 2
Rser 1 3 0.11
Lser 2 4 8.10054347E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885382207011_1nF
*******
.subckt 1206_885382208001_2.2uF 1 2
Rser 1 3 0.011
Lser 2 4 0.0000000011
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885382208001_2.2uF
*******
.subckt 1206_885382208002_10nF 1 2
Rser 1 3 0.131552570055
Lser 2 4 1.072395374E-09
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885382208002_10nF
*******
.subckt 1206_885382208003_100nF 1 2
Rser 1 3 0.0807702333746
Lser 2 4 1.078982226E-09
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885382208003_100nF
*******
.subckt 1206_885382208004_470nF 1 2
Rser 1 3 0.017201291525
Lser 2 4 1.1162727E-12
C1 3 4 0.00000047
Rpar 3 4 1000000000
.ends 1206_885382208004_470nF
*******
.subckt 1206_885382208005_1uF 1 2
Rser 1 3 0.0427768621827
Lser 2 4 1.145259282E-12
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885382208005_1uF
*******
.subckt 1206_885382208006_100nF 1 2
Rser 1 3 0.0371158193445
Lser 2 4 1.097090305E-12
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1206_885382208006_100nF
*******
.subckt 1206_885382208007_100nF 1 2
Rser 1 3 0.03
Lser 2 4 1.025275106E-09
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1206_885382208007_100nF
*******
.subckt 1206_885382208008_270pF 1 2
Rser 1 3 0.00165
Lser 2 4 0.0000000008
C1 3 4 0.00000000027
Rpar 3 4 10000000000
.ends 1206_885382208008_270pF
*******
.subckt 1206_885382208009_10nF 1 2
Rser 1 3 0.0679539884277
Lser 2 4 9.89197769E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885382208009_10nF
*******
.subckt 1206_885382208010_22nF 1 2
Rser 1 3 0.06
Lser 2 4 9.80217377E-10
C1 3 4 0.000000022
Rpar 3 4 4500000000
.ends 1206_885382208010_22nF
*******
.subckt 1206_885382208011_33nF 1 2
Rser 1 3 0.055
Lser 2 4 9.60150263E-10
C1 3 4 0.000000033
Rpar 3 4 3000000000
.ends 1206_885382208011_33nF
*******
.subckt 1206_885382208012_4.7nF 1 2
Rser 1 3 0.11
Lser 2 4 1.00582564E-12
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885382208012_4.7nF
*******
.subckt 1206_885382208013_470pF 1 2
Rser 1 3 0.08
Lser 2 4 8.45206602E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885382208013_470pF
*******
.subckt 1206_885382208014_680pF 1 2
Rser 1 3 0.15
Lser 2 4 8.19920208E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885382208014_680pF
*******
.subckt 1210_885382209001_33nF 1 2
Rser 1 3 0.0375
Lser 2 4 0.000000001
C1 3 4 0.000000033
Rpar 3 4 3000000000
.ends 1210_885382209001_33nF
*******
.subckt 1210_885382209002_2.2uF 1 2
Rser 1 3 0.008
Lser 2 4 0.0000000009
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 1210_885382209002_2.2uF
*******
.subckt 1812_885382211002_100nF 1 2
Rser 1 3 0.0275
Lser 2 4 0.0000000013
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1812_885382211002_100nF
*******
