**************************************************
* Manufacturer:          Würth Elektronik
* Kinds:                 Aluminum Hybrid Polymer Capacitors
* Matchcode:             WCAP-HSAH
* Library Type:          LTspice
* Version:               rev21a
* Created/modified by:   Ella
* Date and Time:         4/26/2023
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************
.subckt 875585344001_100uF 1 2
Rser 1 3 0.024
Lser 2 4 0.00000000275
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 875585344001_100uF
*******
.subckt 875585344003_150uF 1 2
Rser 1 3 0.0189
Lser 2 4 0.00000000275
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 875585344003_150uF
*******
.subckt 875585544002_56uF 1 2
Rser 1 3 0.027
Lser 2 4 0.00000000285
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 875585544002_56uF
*******
.subckt 875585744002_22uF 1 2
Rser 1 3 0.0196
Lser 2 4 0.0000000027
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 875585744002_22uF
*******
.subckt 875585844001_10uF 1 2
Rser 1 3 0.0121
Lser 2 4 0.0000000028
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 875585844001_10uF
*******
.subckt 875585345004_220uF 1 2
Rser 1 3 0.013
Lser 2 4 0.0000000031
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 875585345004_220uF
*******
.subckt 875585545003_100uF 1 2
Rser 1 3 0.014
Lser 2 4 0.0000000031
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 875585545003_100uF
*******
.subckt 875585745003_33uF 1 2
Rser 1 3 0.0145
Lser 2 4 0.000000003
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 875585745003_33uF
*******
.subckt 875585845002_22uF 1 2
Rser 1 3 0.0117
Lser 2 4 0.0000000028
C1 3 4 0.000022
Rpar 3 4 4532374.10071942
.ends 875585845002_22uF
*******
.subckt 875585553004_220uF 1 2
Rser 1 3 0.008
Lser 2 4 0.0000000032
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 875585553004_220uF
*******
.subckt 875585753005_68uF 1 2
Rser 1 3 0.0075
Lser 2 4 0.0000000031
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 875585753005_68uF
*******
.subckt 875585853003_33uF 1 2
Rser 1 3 0.00695
Lser 2 4 0.0000000029
C1 3 4 0.000033
Rpar 3 4 3028846.15384615
.ends 875585853003_33uF
*******
.subckt 875585853004_47uF 1 2
Rser 1 3 0.00715
Lser 2 4 0.0000000031
C1 3 4 0.000047
Rpar 3 4 2128378.37837838
.ends 875585853004_47uF
*******
.subckt 875585357006_330uF 1 2
Rser 1 3 0.0082
Lser 2 4 0.0000000045
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 875585357006_330uF
*******
.subckt 875585357008_470uF 1 2
Rser 1 3 0.0074
Lser 2 4 0.0000000044
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 875585357008_470uF
*******
.subckt 875585357010_560uF 1 2
Rser 1 3 0.0068
Lser 2 4 0.0000000028
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 875585357010_560uF
*******
.subckt 875585557006_330uF 1 2
Rser 1 3 0.0085
Lser 2 4 0.0000000037
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 875585557006_330uF
*******
.subckt 875585757004_56uF 1 2
Rser 1 3 0.0057
Lser 2 4 0.0000000045
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 875585757004_56uF
*******
.subckt 875585757007_100uF 1 2
Rser 1 3 0.0093
Lser 2 4 0.0000000046
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 875585757007_100uF
*******
.subckt 875585857006_56uF 1 2
Rser 1 3 0.0058
Lser 2 4 0.0000000046
C1 3 4 0.000056
Rpar 3 4 1784702.54957507
.ends 875585857006_56uF
*******
.subckt 875585857007_68uF 1 2
Rser 1 3 0.008
Lser 2 4 0.000000004
C1 3 4 0.000068
Rpar 3 4 1471962.61682243
.ends 875585857007_68uF
*******
.subckt 875585957003_22uF 1 2
Rser 1 3 0.0076
Lser 2 4 0.0000000045
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 875585957003_22uF
*******
.subckt 875585361011_820uF 1 2
Rser 1 3 0.0057
Lser 2 4 0.0000000047
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 875585361011_820uF
*******
.subckt 875585561007_470uF 1 2
Rser 1 3 0.006
Lser 2 4 0.0000000037
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 875585561007_470uF
*******
.subckt 875585961005_33uF 1 2
Rser 1 3 0.0084
Lser 2 4 0.0000000041
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 875585961005_33uF
*******
