**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Radial Leaded Wire Wound Inductor
* Matchcode:              WE-TI
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Ella
* Date and Time:          11/9/2022
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 1014_7447480680_68u 1 2
Rp 1 2 67430
Cp 1 2 10.79p
Rs 1 N3 0.063
L1 N3 2 68u
.ends 1014_7447480680_68u
*******
.subckt 1014_7447480101_100u 1 2
Rp 1 2 131910
Cp 1 2 15.5p
Rs 1 N3 0.1
L1 N3 2 100u
.ends 1014_7447480101_100u
*******
.subckt 1014_7447480151_150u 1 2
Rp 1 2 138810
Cp 1 2 16.823p
Rs 1 N3 0.16
L1 N3 2 150u
.ends 1014_7447480151_150u
*******
.subckt 1014_7447480221_220u 1 2
Rp 1 2 140800
Cp 1 2 17.1p
Rs 1 N3 0.23
L1 N3 2 220u
.ends 1014_7447480221_220u
*******
.subckt 1014_7447480331_330u 1 2
Rp 1 2 168000
Cp 1 2 17.4p
Rs 1 N3 0.3
L1 N3 2 330u
.ends 1014_7447480331_330u
*******
.subckt 1014_7447480471_470u 1 2
Rp 1 2 187000
Cp 1 2 17.663p
Rs 1 N3 0.47
L1 N3 2 470u
.ends 1014_7447480471_470u
*******
.subckt 1014_7447480561_560u 1 2
Rp 1 2 100000
Cp 1 2 15.1p
Rs 1 N3 0.55
L1 N3 2 560u
.ends 1014_7447480561_560u
*******
.subckt 1014_7447480681_680u 1 2
Rp 1 2 190350
Cp 1 2 17.8p
Rs 1 N3 0.71
L1 N3 2 680u
.ends 1014_7447480681_680u
*******
.subckt 1014_7447480102_1000u 1 2
Rp 1 2 204700
Cp 1 2 19p
Rs 1 N3 1
L1 N3 2 1000u
.ends 1014_7447480102_1000u
*******
.subckt 1014_7447480122_1200u 1 2
Rp 1 2 214210
Cp 1 2 18p
Rs 1 N3 1.1
L1 N3 2 1200u
.ends 1014_7447480122_1200u
*******
.subckt 1014_7447480152_1500u 1 2
Rp 1 2 270490
Cp 1 2 20.2p
Rs 1 N3 1.5
L1 N3 2 1500u
.ends 1014_7447480152_1500u
*******
.subckt 1014_7447480222_2200u 1 2
Rp 1 2 270490
Cp 1 2 20.2p
Rs 1 N3 2.1
L1 N3 2 2200u
.ends 1014_7447480222_2200u
*******
.subckt 1014_7447480332_3300u 1 2
Rp 1 2 290158
Cp 1 2 18.614p
Rs 1 N3 3.2
L1 N3 2 3300u
.ends 1014_7447480332_3300u
*******
.subckt 1014_7447480562_5600u 1 2
Rp 1 2 332000
Cp 1 2 16p
Rs 1 N3 4.9
L1 N3 2 5600u
.ends 1014_7447480562_5600u
*******
.subckt 1014_7447480822_8200u 1 2
Rp 1 2 290158
Cp 1 2 18.614p
Rs 1 N3 7.5
L1 N3 2 8200u
.ends 1014_7447480822_8200u
*******
.subckt 1016_7447221101_100u 1 2
Rp 1 2 90000
Cp 1 2 14.22p
Rs 1 N3 0.085
L1 N3 2 100u
.ends 1016_7447221101_100u
*******
.subckt 1016_7447221221_220u 1 2
Rp 1 2 107000
Cp 1 2 17.64p
Rs 1 N3 0.19
L1 N3 2 220u
.ends 1016_7447221221_220u
*******
.subckt 1016_7447221331_330u 1 2
Rp 1 2 142600
Cp 1 2 17.7p
Rs 1 N3 0.28
L1 N3 2 330u
.ends 1016_7447221331_330u
*******
.subckt 1016_7447221471_470u 1 2
Rp 1 2 146173.4139506
Cp 1 2 17.02p
Rs 1 N3 0.4
L1 N3 2 470u
.ends 1016_7447221471_470u
*******
.subckt 1016_7447221681_680u 1 2
Rp 1 2 162461.2176448
Cp 1 2 18.84p
Rs 1 N3 0.58
L1 N3 2 680u
.ends 1016_7447221681_680u
*******
.subckt 1016_7447221102_1000u 1 2
Rp 1 2 190000
Cp 1 2 20.02p
Rs 1 N3 0.85
L1 N3 2 1000u
.ends 1016_7447221102_1000u
*******
.subckt 1016_7447221222_2200u 1 2
Rp 1 2 220000
Cp 1 2 18.04p
Rs 1 N3 1.85
L1 N3 2 2200u
.ends 1016_7447221222_2200u
*******
.subckt 1016_7447221332_3300u 1 2
Rp 1 2 254000
Cp 1 2 18.12p
Rs 1 N3 2.8
L1 N3 2 3300u
.ends 1016_7447221332_3300u
*******
.subckt 1016_7447221472_4700u 1 2
Rp 1 2 340000
Cp 1 2 19.1p
Rs 1 N3 4
L1 N3 2 4700u
.ends 1016_7447221472_4700u
*******
.subckt 1016_7447221682_6800u 1 2
Rp 1 2 560000
Cp 1 2 19.3p
Rs 1 N3 5.7
L1 N3 2 6800u
.ends 1016_7447221682_6800u
*******
.subckt 1016_7447221103_10000u 1 2
Rp 1 2 610000
Cp 1 2 21p
Rs 1 N3 8.4
L1 N3 2 10000u
.ends 1016_7447221103_10000u
*******
.subckt 1018_7447231101_100u 1 2
Rp 1 2 100400
Cp 1 2 17.24p
Rs 1 N3 0.075
L1 N3 2 100u
.ends 1018_7447231101_100u
*******
.subckt 1018_7447231221_220u 1 2
Rp 1 2 119000
Cp 1 2 21.96p
Rs 1 N3 0.17
L1 N3 2 220u
.ends 1018_7447231221_220u
*******
.subckt 1018_7447231331_330u 1 2
Rp 1 2 125000
Cp 1 2 20.46p
Rs 1 N3 0.25
L1 N3 2 330u
.ends 1018_7447231331_330u
*******
.subckt 1018_7447231471_470u 1 2
Rp 1 2 147000
Cp 1 2 19.62p
Rs 1 N3 0.36
L1 N3 2 470u
.ends 1018_7447231471_470u
*******
.subckt 1018_7447231681_680u 1 2
Rp 1 2 160000
Cp 1 2 23.5p
Rs 1 N3 0.51
L1 N3 2 680u
.ends 1018_7447231681_680u
*******
.subckt 1018_7447231102_1000u 1 2
Rp 1 2 180280.882332
Cp 1 2 21.68p
Rs 1 N3 0.75
L1 N3 2 1000u
.ends 1018_7447231102_1000u
*******
.subckt 1018_7447231222_2200u 1 2
Rp 1 2 213000
Cp 1 2 20.96p
Rs 1 N3 1.65
L1 N3 2 2200u
.ends 1018_7447231222_2200u
*******
.subckt 1018_7447231332_3300u 1 2
Rp 1 2 259323.969099
Cp 1 2 22.72p
Rs 1 N3 2.45
L1 N3 2 3300u
.ends 1018_7447231332_3300u
*******
.subckt 1018_7447231472_4700u 1 2
Rp 1 2 376000
Cp 1 2 22.78p
Rs 1 N3 3.5
L1 N3 2 4700u
.ends 1018_7447231472_4700u
*******
.subckt 1018_7447231682_6800u 1 2
Rp 1 2 540416.2518812
Cp 1 2 24.3p
Rs 1 N3 5
L1 N3 2 6800u
.ends 1018_7447231682_6800u
*******
.subckt 1018_7447231103_10000u 1 2
Rp 1 2 802741.9933612
Cp 1 2 22.72p
Rs 1 N3 7.4
L1 N3 2 10000u
.ends 1018_7447231103_10000u
*******
.subckt 5075_7447462010_1u 1 2
Rp 1 2 3900
Cp 1 2 1.41p
Rs 1 N3 0.006
L1 N3 2 1u
.ends 5075_7447462010_1u
*******
.subckt 5075_7447462022_2.2u 1 2
Rp 1 2 6700
Cp 1 2 3.06p
Rs 1 N3 0.01
L1 N3 2 2.2u
.ends 5075_7447462022_2.2u
*******
.subckt 5075_7447462033_3.3u 1 2
Rp 1 2 8500
Cp 1 2 3.74p
Rs 1 N3 0.016
L1 N3 2 3.3u
.ends 5075_7447462033_3.3u
*******
.subckt 5075_7447462047_4.7u 1 2
Rp 1 2 10340
Cp 1 2 4.35p
Rs 1 N3 0.019
L1 N3 2 4.7u
.ends 5075_7447462047_4.7u
*******
.subckt 5075_7447462068_6.8u 1 2
Rp 1 2 16020
Cp 1 2 3.78p
Rs 1 N3 0.027
L1 N3 2 6.8u
.ends 5075_7447462068_6.8u
*******
.subckt 5075_7447462100_10u 1 2
Rp 1 2 19570
Cp 1 2 3.53p
Rs 1 N3 0.055
L1 N3 2 10u
.ends 5075_7447462100_10u
*******
.subckt 5075_7447462220_22u 1 2
Rp 1 2 36370
Cp 1 2 5.24p
Rs 1 N3 0.102
L1 N3 2 22u
.ends 5075_7447462220_22u
*******
.subckt 5075_7447462330_33u 1 2
Rp 1 2 49290
Cp 1 2 4.16p
Rs 1 N3 0.153
L1 N3 2 33u
.ends 5075_7447462330_33u
*******
.subckt 5075_7447462470_47u 1 2
Rp 1 2 90960
Cp 1 2 5.43p
Rs 1 N3 0.22
L1 N3 2 47u
.ends 5075_7447462470_47u
*******
.subckt 5075_7447462680_68u 1 2
Rp 1 2 109656
Cp 1 2 6.617p
Rs 1 N3 0.34
L1 N3 2 68u
.ends 5075_7447462680_68u
*******
.subckt 5075_7447462820_82u 1 2
Rp 1 2 63700
Cp 1 2 5.82p
Rs 1 N3 0.39
L1 N3 2 82u
.ends 5075_7447462820_82u
*******
.subckt 5075_7447462101_100u 1 2
Rp 1 2 116350
Cp 1 2 5.47p
Rs 1 N3 0.45
L1 N3 2 100u
.ends 5075_7447462101_100u
*******
.subckt 5075_7447462221_220u 1 2
Rp 1 2 141270
Cp 1 2 8.76p
Rs 1 N3 0.96
L1 N3 2 220u
.ends 5075_7447462221_220u
*******
.subckt 5075_7447462471_470u 1 2
Rp 1 2 162830
Cp 1 2 7.31p
Rs 1 N3 1.58
L1 N3 2 470u
.ends 5075_7447462471_470u
*******
.subckt 5075_7447462681_680u 1 2
Rp 1 2 261612
Cp 1 2 6.983p
Rs 1 N3 3.1
L1 N3 2 680u
.ends 5075_7447462681_680u
*******
.subckt 5075_7447462102_1000u 1 2
Rp 1 2 235800
Cp 1 2 8.48p
Rs 1 N3 4.38
L1 N3 2 1000u
.ends 5075_7447462102_1000u
*******
.subckt 5075_7447462152_1500u 1 2
Rp 1 2 582140
Cp 1 2 9.7p
Rs 1 N3 6.54
L1 N3 2 1500u
.ends 5075_7447462152_1500u
*******
.subckt 5075_7447462222_2200u 1 2
Rp 1 2 611898
Cp 1 2 9.38p
Rs 1 N3 9.8
L1 N3 2 2200u
.ends 5075_7447462222_2200u
*******
.subckt 6065_744779068_6.8u 1 2
Rp 1 2 16190
Cp 1 2 2.94p
Rs 1 N3 0.027
L1 N3 2 6.8u
.ends 6065_744779068_6.8u
*******
.subckt 6065_744779100_10u 1 2
Rp 1 2 19660
Cp 1 2 3.53p
Rs 1 N3 0.0386
L1 N3 2 10u
.ends 6065_744779100_10u
*******
.subckt 6065_7447790470_47u 1 2
Rp 1 2 61680
Cp 1 2 5.66p
Rs 1 N3 0.135
L1 N3 2 47u
.ends 6065_7447790470_47u
*******
.subckt 6065_744779168_68u 1 2
Rp 1 2 65000
Cp 1 2 4.2p
Rs 1 N3 0.22
L1 N3 2 68u
.ends 6065_744779168_68u
*******
.subckt 6065_7447790221_220u 1 2
Rp 1 2 193000
Cp 1 2 5.81p
Rs 1 N3 0.64
L1 N3 2 220u
.ends 6065_7447790221_220u
*******
.subckt 8012_7447452100_10u 1 2
Rp 1 2 13360
Cp 1 2 7.93p
Rs 1 N3 0.015
L1 N3 2 10u
.ends 8012_7447452100_10u
*******
.subckt 8012_7447452101_100u 1 2
Rp 1 2 113550
Cp 1 2 12.24p
Rs 1 N3 0.13
L1 N3 2 100u
.ends 8012_7447452101_100u
*******
.subckt 8012_7447452221_220u 1 2
Rp 1 2 151910
Cp 1 2 13.361p
Rs 1 N3 0.27
L1 N3 2 220u
.ends 8012_7447452221_220u
*******
.subckt 8012_7447452331_330u 1 2
Rp 1 2 156320
Cp 1 2 14.007p
Rs 1 N3 0.42
L1 N3 2 330u
.ends 8012_7447452331_330u
*******
.subckt 8012_7447452391_390u 1 2
Rp 1 2 204810
Cp 1 2 13.933p
Rs 1 N3 0.47
L1 N3 2 390u
.ends 8012_7447452391_390u
*******
.subckt 8012_7447452561_560u 1 2
Rp 1 2 199096
Cp 1 2 13.363p
Rs 1 N3 0.69
L1 N3 2 560u
.ends 8012_7447452561_560u
*******
.subckt 8012_7447452821_820u 1 2
Rp 1 2 251962
Cp 1 2 12.755p
Rs 1 N3 1
L1 N3 2 820u
.ends 8012_7447452821_820u
*******
.subckt 8012_7447452102_1000u 1 2
Rp 1 2 206258
Cp 1 2 12.713p
Rs 1 N3 1.27
L1 N3 2 1000u
.ends 8012_7447452102_1000u
*******
.subckt 8012_7447452152_1500u 1 2
Rp 1 2 286306
Cp 1 2 15.581p
Rs 1 N3 1.75
L1 N3 2 1500u
.ends 8012_7447452152_1500u
*******
.subckt 8012_7447452222_2200u 1 2
Rp 1 2 299390
Cp 1 2 12.654p
Rs 1 N3 2.4
L1 N3 2 2200u
.ends 8012_7447452222_2200u
*******
.subckt 8012_7447452392_3900u 1 2
Rp 1 2 568880
Cp 1 2 14.285p
Rs 1 N3 4.55
L1 N3 2 3900u
.ends 8012_7447452392_3900u
*******
.subckt 8012_7447452472_4700u 1 2
Rp 1 2 695000
Cp 1 2 14.368p
Rs 1 N3 6.1
L1 N3 2 4700u
.ends 8012_7447452472_4700u
*******
.subckt 8012_7447452103_10000u 1 2
Rp 1 2 500000
Cp 1 2 13p
Rs 1 N3 13
L1 N3 2 10000u
.ends 8012_7447452103_10000u
*******
.subckt 8012_7447452683_68000u 1 2
Rp 1 2 709600
Cp 1 2 15.406p
Rs 1 N3 90
L1 N3 2 68000u
.ends 8012_7447452683_68000u
*******
.subckt 8012_7447450103_10000u 1 2
Rp 1 2 447280
Cp 1 2 12.987p
Rs 1 N3 13
L1 N3 2 10000u
.ends 8012_7447450103_10000u
*******
.subckt 8012B_744743101_100u 1 2
Rp 1 2 89830
Cp 1 2 10.34p
Rs 1 N3 0.25
L1 N3 2 100u
.ends 8012B_744743101_100u
*******
.subckt 8012B_744743221_220u 1 2
Rp 1 2 129470
Cp 1 2 9.45p
Rs 1 N3 0.47
L1 N3 2 220u
.ends 8012B_744743221_220u
*******
.subckt 8012B_744743331_330u 1 2
Rp 1 2 141390
Cp 1 2 10.41p
Rs 1 N3 0.97
L1 N3 2 330u
.ends 8012B_744743331_330u
*******
.subckt 8012B_744743471_470u 1 2
Rp 1 2 156110
Cp 1 2 12.85p
Rs 1 N3 1.13
L1 N3 2 470u
.ends 8012B_744743471_470u
*******
.subckt 8012B_744743102_1000u 1 2
Rp 1 2 165950
Cp 1 2 13.4p
Rs 1 N3 2.24
L1 N3 2 1000u
.ends 8012B_744743102_1000u
*******
.subckt 8055_744741101_100u 1 2
Rp 1 2 78440
Cp 1 2 3.48p
Rs 1 N3 0.42
L1 N3 2 100u
.ends 8055_744741101_100u
*******
.subckt 8055_744741221_220u 1 2
Rp 1 2 103200
Cp 1 2 4.52p
Rs 1 N3 0.97
L1 N3 2 220u
.ends 8055_744741221_220u
*******
.subckt 8055_7447412331_330u 1 2
Rp 1 2 115850
Cp 1 2 4.82p
Rs 1 N3 1.25
L1 N3 2 330u
.ends 8055_7447412331_330u
*******
.subckt 8055_744741471_470u 1 2
Rp 1 2 158980
Cp 1 2 4.95p
Rs 1 N3 2.12
L1 N3 2 470u
.ends 8055_744741471_470u
*******
.subckt 8055_7447412681_680u 1 2
Rp 1 2 160310
Cp 1 2 5p
Rs 1 N3 2.62
L1 N3 2 680u
.ends 8055_7447412681_680u
*******
.subckt 8055_744741102_1000u 1 2
Rp 1 2 220000
Cp 1 2 5.685p
Rs 1 N3 4.49
L1 N3 2 1000u
.ends 8055_744741102_1000u
*******
.subckt 8055_744741222_2200u 1 2
Rp 1 2 225450
Cp 1 2 5.88p
Rs 1 N3 9.13
L1 N3 2 2200u
.ends 8055_744741222_2200u
*******
.subckt 8055_744741472_4700u 1 2
Rp 1 2 500000
Cp 1 2 6.12p
Rs 1 N3 21.18
L1 N3 2 4700u
.ends 8055_744741472_4700u
*******
.subckt 8075_744732015_1.5u 1 2
Rp 1 2 4350
Cp 1 2 1.45p
Rs 1 N3 0.007
L1 N3 2 1.5u
.ends 8075_744732015_1.5u
*******
.subckt 8075_744732100_10u 1 2
Rp 1 2 21050
Cp 1 2 4.24p
Rs 1 N3 0.027
L1 N3 2 10u
.ends 8075_744732100_10u
*******
.subckt 8075_744732470_47u 1 2
Rp 1 2 48547
Cp 1 2 8.51p
Rs 1 N3 0.114
L1 N3 2 47u
.ends 8075_744732470_47u
*******
.subckt 8075_744732121_120u 1 2
Rp 1 2 82430
Cp 1 2 6.29p
Rs 1 N3 0.34
L1 N3 2 120u
.ends 8075_744732121_120u
*******
.subckt 8075_744732221_220u 1 2
Rp 1 2 162670
Cp 1 2 5.83p
Rs 1 N3 0.59
L1 N3 2 220u
.ends 8075_744732221_220u
*******
.subckt 8075_744732331_330u 1 2
Rp 1 2 199060
Cp 1 2 5.38p
Rs 1 N3 0.94
L1 N3 2 330u
.ends 8075_744732331_330u
*******
.subckt 8075_744732471_470u 1 2
Rp 1 2 273530
Cp 1 2 6.69p
Rs 1 N3 1.44
L1 N3 2 470u
.ends 8075_744732471_470u
*******
.subckt 8075_744732681_680u 1 2
Rp 1 2 283430
Cp 1 2 7.94p
Rs 1 N3 1.79
L1 N3 2 680u
.ends 8075_744732681_680u
*******
.subckt 8075_744732102_1000u 1 2
Rp 1 2 314850
Cp 1 2 7.73p
Rs 1 N3 2.8
L1 N3 2 1000u
.ends 8075_744732102_1000u
*******
.subckt 8075_744732152_1500u 1 2
Rp 1 2 500000
Cp 1 2 4.5p
Rs 1 N3 4.25
L1 N3 2 1500u
.ends 8075_744732152_1500u
*******
.subckt 8075_744730392_3900u 1 2
Rp 1 2 534741.4
Cp 1 2 4.6339p
Rs 1 N3 9.5
L1 N3 2 3900u
.ends 8075_744730392_3900u
*******
.subckt 8075_7447721047_4700u 1 2
Rp 1 2 358840
Cp 1 2 6.93p
Rs 1 N3 10.98
L1 N3 2 4700u
.ends 8075_7447721047_4700u
*******
.subckt 8075_744732153_15000u 1 2
Rp 1 2 1300000
Cp 1 2 8p
Rs 1 N3 50
L1 N3 2 15000u
.ends 8075_744732153_15000u
*******
.subckt 8095_7447720010_1u 1 2
Rp 1 2 3241
Cp 1 2 0.873729p
Rs 1 N3 0.009
L1 N3 2 0.773822u
.ends 8095_7447720010_1u
*******
.subckt 8095_7447720022_2.2u 1 2
Rp 1 2 6702
Cp 1 2 0.855743p
Rs 1 N3 0.013
L1 N3 2 1.946u
.ends 8095_7447720022_2.2u
*******
.subckt 8095_7447720033_3.3u 1 2
Rp 1 2 10043
Cp 1 2 0.882163p
Rs 1 N3 0.016
L1 N3 2 3.01u
.ends 8095_7447720033_3.3u
*******
.subckt 8095_7447720047_4.7u 1 2
Rp 1 2 13.136
Cp 1 2 1.153p
Rs 1 N3 0.019
L1 N3 2 4.406u
.ends 8095_7447720047_4.7u
*******
.subckt 8095_7447720068_6.8u 1 2
Rp 1 2 10285
Cp 1 2 2.68p
Rs 1 N3 0.024
L1 N3 2 6.988u
.ends 8095_7447720068_6.8u
*******
.subckt 8095_7447720100_10u 1 2
Rp 1 2 11820
Cp 1 2 7.309p
Rs 1 N3 0.03
L1 N3 2 9.913u
.ends 8095_7447720100_10u
*******
.subckt 8095_7447720150_15u 1 2
Rp 1 2 18894
Cp 1 2 6.393p
Rs 1 N3 0.038
L1 N3 2 15.024u
.ends 8095_7447720150_15u
*******
.subckt 8095_7447720180_18u 1 2
Rp 1 2 19905
Cp 1 2 5.974p
Rs 1 N3 0.042
L1 N3 2 18.111u
.ends 8095_7447720180_18u
*******
.subckt 8095_7447720200_20u 1 2
Rp 1 2 24975
Cp 1 2 5.532p
Rs 1 N3 0.044
L1 N3 2 19.302u
.ends 8095_7447720200_20u
*******
.subckt 8095_7447720220_22u 1 2
Rp 1 2 19554
Cp 1 2 7.128p
Rs 1 N3 0.046
L1 N3 2 20.467u
.ends 8095_7447720220_22u
*******
.subckt 8095_7447720330_33u 1 2
Rp 1 2 28146
Cp 1 2 6.327p
Rs 1 N3 0.059
L1 N3 2 30.792u
.ends 8095_7447720330_33u
*******
.subckt 8095_7447720390_39u 1 2
Rp 1 2 31820
Cp 1 2 6.363p
Rs 1 N3 0.07
L1 N3 2 37.353u
.ends 8095_7447720390_39u
*******
.subckt 8095_7447720470_47u 1 2
Rp 1 2 43543
Cp 1 2 6.501p
Rs 1 N3 0.089
L1 N3 2 46.318u
.ends 8095_7447720470_47u
*******
.subckt 8095_7447720560_56u 1 2
Rp 1 2 41474
Cp 1 2 7.011p
Rs 1 N3 0.1
L1 N3 2 52.525u
.ends 8095_7447720560_56u
*******
.subckt 8095_7447720680_68u 1 2
Rp 1 2 44794
Cp 1 2 8.66p
Rs 1 N3 0.124
L1 N3 2 64.373u
.ends 8095_7447720680_68u
*******
.subckt 8095_7447720820_82u 1 2
Rp 1 2 52955
Cp 1 2 8.192p
Rs 1 N3 0.154
L1 N3 2 80.317u
.ends 8095_7447720820_82u
*******
.subckt 8095_7447720101_100u 1 2
Rp 1 2 78404
Cp 1 2 6.957p
Rs 1 N3 0.198
L1 N3 2 97.702u
.ends 8095_7447720101_100u
*******
.subckt 8095_7447720121_120u 1 2
Rp 1 2 69934
Cp 1 2 7.531p
Rs 1 N3 0.223
L1 N3 2 113.151u
.ends 8095_7447720121_120u
*******
.subckt 8095_7447720151_150u 1 2
Rp 1 2 85014
Cp 1 2 8.411p
Rs 1 N3 0.283
L1 N3 2 147.802u
.ends 8095_7447720151_150u
*******
.subckt 8095_7447720181_180u 1 2
Rp 1 2 80820
Cp 1 2 9.507p
Rs 1 N3 0.35
L1 N3 2 184.96u
.ends 8095_7447720181_180u
*******
.subckt 8095_7447720221_220u 1 2
Rp 1 2 96670
Cp 1 2 8.194p
Rs 1 N3 0.389
L1 N3 2 211.021u
.ends 8095_7447720221_220u
*******
.subckt 8095_7447720331_330u 1 2
Rp 1 2 128923
Cp 1 2 7.838p
Rs 1 N3 0.587
L1 N3 2 322.954u
.ends 8095_7447720331_330u
*******
.subckt 8095_7447720471_470u 1 2
Rp 1 2 129153
Cp 1 2 9.486p
Rs 1 N3 0.883
L1 N3 2 462.051u
.ends 8095_7447720471_470u
*******
.subckt 8095_7447720561_560u 1 2
Rp 1 2 161978
Cp 1 2 8.314p
Rs 1 N3 1.02
L1 N3 2 551.143u
.ends 8095_7447720561_560u
*******
.subckt 8095_7447720681_680u 1 2
Rp 1 2 177759
Cp 1 2 8.457p
Rs 1 N3 1.29
L1 N3 2 664.793u
.ends 8095_7447720681_680u
*******
.subckt 8095_7447720821_820u 1 2
Rp 1 2 167440
Cp 1 2 7.888p
Rs 1 N3 1.41
L1 N3 2 775.226u
.ends 8095_7447720821_820u
*******
.subckt 8095_7447720901_900u 1 2
Rp 1 2 205905
Cp 1 2 8.509p
Rs 1 N3 1.68
L1 N3 2 862.244u
.ends 8095_7447720901_900u
*******
.subckt 8095_7447720102_1000u 1 2
Rp 1 2 206222
Cp 1 2 8.97p
Rs 1 N3 1.89
L1 N3 2 1001u
.ends 8095_7447720102_1000u
*******
.subckt 8095_7447720122_1200u 1 2
Rp 1 2 195247
Cp 1 2 8.535p
Rs 1 N3 2.14
L1 N3 2 1182u
.ends 8095_7447720122_1200u
*******
.subckt 8095_7447720152_1500u 1 2
Rp 1 2 207270
Cp 1 2 8.972p
Rs 1 N3 2.67
L1 N3 2 1460u
.ends 8095_7447720152_1500u
*******
.subckt 8095_7447720182_1800u 1 2
Rp 1 2 293012
Cp 1 2 8.157p
Rs 1 N3 3.68
L1 N3 2 1757u
.ends 8095_7447720182_1800u
*******
.subckt 8095_7447720222_2200u 1 2
Rp 1 2 288136
Cp 1 2 8.535p
Rs 1 N3 4.16
L1 N3 2 2152u
.ends 8095_7447720222_2200u
*******
.subckt 8095_7447720332_3300u 1 2
Rp 1 2 303912
Cp 1 2 8.123p
Rs 1 N3 6.53
L1 N3 2 3237u
.ends 8095_7447720332_3300u
*******
.subckt 8095_7447720392_3900u 1 2
Rp 1 2 472730
Cp 1 2 8.446p
Rs 1 N3 7.34
L1 N3 2 3847u
.ends 8095_7447720392_3900u
*******
.subckt 8095_7447720472_4700u 1 2
Rp 1 2 476334
Cp 1 2 7.879p
Rs 1 N3 8.33
L1 N3 2 4636u
.ends 8095_7447720472_4700u
*******
.subckt 8095_7447720702_7000u 1 2
Rp 1 2 472208
Cp 1 2 7.297p
Rs 1 N3 13.3
L1 N3 2 6767u
.ends 8095_7447720702_7000u
*******
.subckt 8095_7447720103_10000u 1 2
Rp 1 2 567589
Cp 1 2 9.307p
Rs 1 N3 19.52
L1 N3 2 9858u
.ends 8095_7447720103_10000u
*******
.subckt 8095_7447720223_22000u 1 2
Rp 1 2 958933
Cp 1 2 7.859p
Rs 1 N3 43.23
L1 N3 2 21899u
.ends 8095_7447720223_22000u
*******
.subckt 8095_7447722363_36000u 1 2
Rp 1 2 1740000
Cp 1 2 10.671p
Rs 1 N3 69.7
L1 N3 2 35500u
.ends 8095_7447722363_36000u
*******
.subckt 8095_7447722473_47000u 1 2
Rp 1 2 1630000
Cp 1 2 10.685p
Rs 1 N3 90.8
L1 N3 2 47493u
.ends 8095_7447722473_47000u
*******
