**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Current Sense Transformer
* Matchcode:              WE-CST 
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Toby      
* Date and Time:          2022-09-13
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************	
.subckt	749252020		3  4  1  2		
.param RxLkg=43.56ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	48.8uH	Rser=290mohm	
K Lpri1    Lsec1        1					
.param Cprm1=1080pf					
.param Rdmp1=531.42ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					
	

.subckt	749252030		3  4  1  2		
.param RxLkg=29.04ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	109.8uH	Rser=660mohm	
K Lpri1    Lsec1        1					
.param Cprm1=2430pf					
.param Rdmp1=354.28ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					
	

.subckt	749252040		3  4  1  2		
.param RxLkg=21.78ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	195.2uH	Rser=1030mohm	
K Lpri1    Lsec1        1					
.param Cprm1=4320pf					
.param Rdmp1=265.71ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					
	

.subckt	749252050		3  4  1  2		
.param RxLkg=17.42ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	305uH	Rser=1660mohm	
K Lpri1    Lsec1        1					
.param Cprm1=6750pf					
.param Rdmp1=212.57ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					
		

.subckt	749252060		3  4  1  2		
.param RxLkg=14.52ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	439.2uH	Rser=2530mohm	
K Lpri1    Lsec1        1					
.param Cprm1=9720pf					
.param Rdmp1=177.14ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					
		

.subckt	749252070		3  4  1  2		
.param RxLkg=12.45ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	597.8uH	Rser=3730mohm	
K Lpri1    Lsec1        1					
.param Cprm1=13230pf					
.param Rdmp1=151.83ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					
		

.subckt	749252100		3  4  1  2		
.param RxLkg=8.71ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	1220uH	Rser=7060mohm	
K Lpri1    Lsec1        1					
.param Cprm1=27000pf					
.param Rdmp1=106.28ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					
		

.subckt	749252125		3  4  1  2		
.param RxLkg=6.97ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	1906.25uH	Rser=10440mohm	
K Lpri1    Lsec1        1					
.param Cprm1=42187pf					
.param Rdmp1=85.03ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					

.subckt	749252150		3  4  1  2		
.param RxLkg=5.81ohm					
.param Leakage=0.01uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.001mohm	
Lpri1	3a	4	0.112uH	Rser=2.3mohm	
Lsec1	1	2	2745uH	Rser=15530mohm	
K Lpri1    Lsec1        1					
.param Cprm1=60750pf					
.param Rdmp1=70.86ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	1	0	20meg		
Rg19	2	0	20meg		
.ends					


.subckt	749251020		8  7  1  3		
.param RxLkg=8.42ohm					
.param Leakage=0.0035uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.297uH	Rser=0.55mohm	
Lsec1	1	3	120uH	Rser=160mohm	
K Lpri1    Lsec1        1					
.param Cprm1=1440pf					
.param Rdmp1=721.69ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					


.subckt	749251030		8  7  1  3		
.param RxLkg=5.3ohm					
.param Leakage=0.0035uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.297uH	Rser=0.55mohm	
Lsec1	1	3	270uH	Rser=396mohm	
K Lpri1    Lsec1        1					
.param Cprm1=3630pf					
.param Rdmp1=454.55ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					

.subckt	749251040		8  7  1  3		
.param RxLkg=3.32ohm					
.param Leakage=0.0035uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.297uH	Rser=0.55mohm	
Lsec1	1	3	480uH	Rser=683mohm	
K Lpri1    Lsec1        1					
.param Cprm1=9235pf					
.param Rdmp1=284.98ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					

.subckt	749251050		8  7  1  3		
.param RxLkg=2.37ohm					
.param Leakage=0.0035uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.297uH	Rser=0.55mohm	
Lsec1	1	3	750uH	Rser=1030mohm	
K Lpri1    Lsec1        1					
.param Cprm1=18170pf					
.param Rdmp1=203.17ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					


.subckt	749251060		8  7  1  3		
.param RxLkg=2.05ohm					
.param Leakage=0.0035uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.297uH	Rser=0.55mohm	
Lsec1	1	3	1080uH	Rser=1492mohm	
K Lpri1    Lsec1        1					
.param Cprm1=24400pf					
.param Rdmp1=175.32ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					


.subckt	749251070		8  7  1  3		
.param RxLkg=1.68ohm					
.param Leakage=0.0035uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.297uH	Rser=0.55mohm	
Lsec1	1	3	1470uH	Rser=1772mohm	
K Lpri1    Lsec1        1					
.param Cprm1=36201pf					
.param Rdmp1=143.94ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					
	

.subckt	749251100		8  7  1  3		
.param RxLkg=1.18ohm					
.param Leakage=0.0035uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.297uH	Rser=0.55mohm	
Lsec1	1	3	3000uH	Rser=3886mohm	
K Lpri1    Lsec1        1					
.param Cprm1=73540pf					
.param Rdmp1=100.99ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					

.subckt	749251125		8  7  1  3		
.param RxLkg=0.96ohm					
.param Leakage=0.0035uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.297uH	Rser=0.55mohm	
Lsec1	1	3	4687.5uH	Rser=4894mohm	
K Lpri1    Lsec1        1					
.param Cprm1=111406pf					
.param Rdmp1=82.05ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					

.subckt	749251150		8  7  1  3		
.param RxLkg=1.71ohm					
.param Leakage=0.009uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.291uH	Rser=0.55mohm	
Lsec1	1	3	6750uH	Rser=8044mohm	
K Lpri1    Lsec1        1					
.param Cprm1=231750pf					
.param Rdmp1=56.89ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					
	

.subckt	749251200		8  7  1  3		
.param RxLkg=1.4ohm					
.param Leakage=0.008uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.292uH	Rser=0.55mohm	
Lsec1	1	3	12000uH	Rser=14180mohm	
K Lpri1    Lsec1        1					
.param Cprm1=271200pf					
.param Rdmp1=52.59ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					


.subckt	749251250		8  7  1  3		
.param RxLkg=0.75ohm					
.param Leakage=0.007uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.001mohm	
Lpri1	8a	7	0.293uH	Rser=0.55mohm	
Lsec1	1	3	18750uH	Rser=19940mohm	
K Lpri1    Lsec1        1					
.param Cprm1=718750pf					
.param Rdmp1=32.3ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg7	7	0	20meg		
Rg11	1	0	20meg		
Rg19	3	0	20meg		
.ends					
	
	
.subckt	7492540020		11  12  2  4		
.param RxLkg=5.37ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	340uH	Rser=33mohm	
K Lpri1    Lsec1        1					
.param Cprm1=5000pf					
.param Rdmp1=651.92ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					
		

.subckt	7492540030		11  12  2  4		
.param RxLkg=2.96ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	765uH	Rser=93mohm	
K Lpri1    Lsec1        1					
.param Cprm1=16500pf					
.param Rdmp1=358.87ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					

.subckt	7492540040		11  12  2  4		
.param RxLkg=2.27ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	1360uH	Rser=130mohm	
K Lpri1    Lsec1        1					
.param Cprm1=28000pf					
.param Rdmp1=275.48ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					
		

.subckt	7492540050		11  12  2  4		
.param RxLkg=1.71ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	2125uH	Rser=202mohm	
K Lpri1    Lsec1        1					
.param Cprm1=49500pf					
.param Rdmp1=207.19ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					
	

.subckt	7492540060		11  12  2  4		
.param RxLkg=1.35ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	3060uH	Rser=305mohm	
K Lpri1    Lsec1        1					
.param Cprm1=79000pf					
.param Rdmp1=164.01ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					
	

.subckt	7492540070		11  12  2  4		
.param RxLkg=1.2ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	4165uH	Rser=367mohm	
K Lpri1    Lsec1        1					
.param Cprm1=100000pf					
.param Rdmp1=145.77ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					
	

.subckt	7492540100		11  12  2  4		
.param RxLkg=0.85ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	8500uH	Rser=805mohm	
K Lpri1    Lsec1        1					
.param Cprm1=200000pf					
.param Rdmp1=103.08ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					

.subckt	7492540150		11  12  2  4		
.param RxLkg=0.58ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	19125uH	Rser=1900mohm	
K Lpri1    Lsec1        1					
.param Cprm1=425000pf					
.param Rdmp1=70.71ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					
	

.subckt	7492540200		11  12  2  4		
.param RxLkg=0.34ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	34000uH	Rser=2630mohm	
K Lpri1    Lsec1        1					
.param Cprm1=1250000pf					
.param Rdmp1=41.23ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					

.subckt	7492540500		11  12  2  4		
.param RxLkg=0.16ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	212500uH	Rser=21200mohm	
K Lpri1    Lsec1        1					
.param Cprm1=5580000pf					
.param Rdmp1=19.51ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					
	

.subckt	7492540750		11  12  2  4		
.param RxLkg=0.1ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	478125uH	Rser=50100mohm	
K Lpri1    Lsec1        1					
.param Cprm1=14200000pf					
.param Rdmp1=12.24ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					

.subckt	7492541000		11  12  2  4		
.param RxLkg=0.08ohm					
.param Leakage=0.007uh					
Rlkg	11	11a	{RxLkg}		
L_Lkg	11	11a	{Leakage}	Rser=0.001mohm	
Lpri1	11a	12	0.843uH	Rser=0.2mohm	
Lsec1	2	4	850000uH	Rser=87640mohm	
K Lpri1    Lsec1        1					
.param Cprm1=21200000pf					
.param Rdmp1=10.01ohm					
Cpri1	11	12	{Cprm1}	Rser=10mohm	
Rdmp1	11	12	{Rdmp1}		
Rg3	11	0	20meg		
Rg7	12	0	20meg		
Rg11	2	0	20meg		
Rg19	4	0	20meg		
.ends					

		