**************************************************
* Manufacturer:           Würth Elektronik 
* Kinds:                  Ferrite SMT Inductor
* Matchcode:              WE-RFI 
* Library Type:           LTspice
* Version:                rev24a
* Created/modified by:    Ella      
* Date and Time:          2024-03-06
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2024 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0402_7447650120_0.02u 1 2
C1 1 N7 13.7521p
L1 1 N1 17.4870n
L2 N1 N2 41.2872p
L3 N2 N3 452.0712p
L4 N3 N4 1.4331n
L5 N4 N5 1.5877n
L6 N5 N6 2.0026n
R1 2 N1 3.9201
R2 2 N2 4.6868
R3 2 N3 1.1576
R4 2 N4 232.2617m
R5 2 N5 50.5841m
R6 2 N6 27.6518m
R7 2 N7 190.4193
R8 2 1 10g
.ends 
*******
.subckt 0402_7447650130_0.03u 1 2
C1 1 N7 74.1373f
L1 1 N1 28.1000n
L2 N1 N2 39.3860p
L3 N2 N3 377.5031p
L4 N3 N4 1.7080n
L5 N4 N5 1.8696n
L6 N5 N6 4.3651n
R1 2 N1 1.8834
R2 2 N2 1.6424
R3 2 N3 1.1069
R4 2 N4 338.3874m
R5 2 N5 61.5372m
R6 2 N6 43.7882m
R7 2 N7 3.7356
R8 2 1 10G
R9 2 1 247.8412
.ends 
*******
.subckt 0402_7447650133_0.033u 1 2
C1 1 N7 43f
L1 1 N1 30n
L2 N1 N2 3.2546p
L3 N2 N3 7.9174p
L4 N3 N4 2.3144n
L5 N4 N5 2.3746n
L6 N5 N6 9.0699n
R1 2 N1 2.4410
R2 2 N2 2.3552
R3 2 N3 2.3004
R4 2 N4 416.0870m
R5 2 N5 67.4299m
R6 2 N6 55.6156m
R7 2 N7 3.7348
R8 2 1 10G
R9 2 1 302.1007
.ends 
*******
.subckt 0402_7447650136_0.036u 1 2
C1 1 N7 46f
L1 1 N1 33n
L2 N1 N2 6.6183p
L3 N2 N3 1.2288n
L4 N3 N4 2.7651n
L5 N4 N5 2.7630n
L6 N5 N6 8.2439n
R1 2 N1 1.8714
R2 2 N2 1.8998
R3 2 N3 1.3853
R4 2 N4 149.8217m
R5 2 N5 95.1510m
R6 2 N6 70.4428m
R7 2 N7 4.0936
R8 2 1 10G
R9 2 1 380
.ends 
*******
.subckt 0402_7447650177_0.077u 1 2
C1 1 N7 40.4951f
L1 1 N1 69.3961n
L2 N1 N2 6.5991p
L3 N2 N3 3.7914n
L4 N3 N4 2.8741n
L5 N4 N5 2.0992n
L6 N5 N6 9.8267n
R1 2 N1 5.8992
R2 2 N2 1.9172
R3 2 N3 6.3978
R4 2 N4 7.0023
R5 2 N5 187.0550m
R6 2 N6 109.6122m
R7 2 N7 9.9867
R8 2 1 10G
R9 2 1 767.8726
.ends 
*******
.subckt 0402_7447650190_0.09u 1 2
C1 1 N7 35.4057f
L1 1 N1 80.0700n
L2 N1 N2 805.6234p
L3 N2 N3 9.5671n
L4 N3 N4 8.0140n
L5 N4 N5 68.0257p
L6 N5 N6 42.7803p
R1 2 N1 8.1400
R2 2 N2 2.4557
R3 2 N3 354.5040m
R4 2 N4 248.0783m
R5 2 N5 408.5573m
R6 2 N6 420.6439m
R7 2 N7 10.3973
R8 2 1 10G
R9 2 1 1.0005k
.ends 
*******
.subckt 0402_7447650210_0.1u 1 2
C1 1 N7 40.6443f
L1 1 N1 88n
L2 N1 N2 1.0040n
L3 N2 N3 8.4138n
L4 N3 N4 8.6302n
L5 N4 N5 1.0012n
L6 N5 N6 676.7281p
R1 2 N1 11.0819
R2 2 N2 4.8111
R3 2 N3 636.7791m
R4 2 N4 875.8463m
R5 2 N5 876.1176m
R6 2 N6 175.3248m
R7 2 N7 10.3669
R8 2 1 10G
R9 2 1 1.1743k
.ends 
*******
.subckt 0402_7447650212_0.12u 1 2
C1 1 N7 30.9067f
L1 1 N1 108.1887n
L2 N1 N2 95.5213p
L3 N2 N3 10.0074n
L4 N3 N4 9.7912n
L5 N4 N5 2.8734n
L6 N5 N6 692.6247p
R1 2 N1 9.4239
R2 2 N2 4.7262
R3 2 N3 781.4822m
R4 2 N4 882.2140m
R5 2 N5 879.2858m
R6 2 N6 205.7003m
R7 2 N7 10.3929
R8 2 1 10G
R9 2 1 1.2062k
.ends 
*******
.subckt 0402_7447650215_0.15u 1 2
C1 1 N7 29.0305f
L1 1 N1 135.0125n
L2 N1 N2 30.3877p
L3 N2 N3 11.5408n
L4 N3 N4 8.4700n
L5 N4 N5 12.5710n
L6 N5 N6 11.2926n
R1 2 N1 7.1528
R2 2 N2 8.1543
R3 2 N3 3.3215
R4 2 N4 255.8154m
R5 2 N5 121.9879m
R6 2 N6 413.4272m
R7 2 N7 10.8114
R8 2 1 10G
R9 2 1 1.9715k
.ends 
*******
.subckt 0402_7447650218_0.18u 1 2
C1 1 N7 23.7055f
L1 1 N1 162.2169n
L2 N1 N2 5.9513p
L3 N2 N3 11.6093n
L4 N3 N4 9.4895n
L5 N4 N5 12.7600n
L6 N5 N6 22.1667n
R1 2 N1 12.0127
R2 2 N2 6.1888
R3 2 N3 2.5800
R4 2 N4 401.8570m
R5 2 N5 315.7505m
R6 2 N6 272.1154m
R7 2 N7 4.0931
R8 2 1 10G
R9 2 1 1.7180k
.ends 
*******
.subckt 0402_7447650222_0.22u 1 2
C1 1 N7 28.5525f
L1 1 N1 197.8283n
L2 N1 N2 45.8140p
L3 N2 N3 10.2070n
L4 N3 N4 16.5065n
L5 N4 N5 19.0510n
L6 N5 N6 42.1733n
R1 2 N1 14.6050
R2 2 N2 13.7443
R3 2 N3 10.0910
R4 2 N4 551.8277m
R5 2 N5 435.0831m
R6 2 N6 691.2797m
R7 2 N7 4.0935
R8 2 1 10G
R9 2 1 2.3240k
.ends 
*******
.subckt 0402_7447650227_0.27u 1 2
C1 1 N7 23.5525f
L1 1 N1 243.8283n
L2 N1 N2 45.8107p
L3 N2 N3 9.0687n
L4 N3 N4 21.7873n
L5 N4 N5 33.9583n
L6 N5 N6 43.6065n
R1 2 N1 14.5358
R2 2 N2 13.6661
R3 2 N3 10.0208
R4 2 N4 636.2071m
R5 2 N5 485.8146m
R6 2 N6 690.2297m
R7 2 N7 4.0935
R8 2 1 10G
R9 2 1 2.7240kA
.ends 
*******
.subckt 0402_7447650233_0.33u 1 2
C1 1 N7 40.5634f
L1 1 N1 287n
L2 N1 N2 7045.5386p
L3 N2 N3 11.6011n
L4 N3 N4 23.2715n
L5 N4 N5 26.7286n
L6 N5 N6 98.2395n
R1 2 N1 78.5804
R2 2 N2 46.7639
R3 2 N3 38.1444
R4 2 N4 2.2482
R5 2 N5 612.3127m
R6 2 N6 221.5058m
R7 2 N7 40.1597
R8 2 1 10G
R9 2 1 4.3021k
.ends 
*******
.subckt 0402_7447650236_0.36u 1 2
C1 1 N7 32.8327f
L1 1 N1 312.8953n
L2 N1 N2 7.1304n
L3 N2 N3 3.3486n
L4 N3 N4 28.8441n
L5 N4 N5 30.8457n
L6 N5 N6 105.8701n
R1 2 N1 78.5104
R2 2 N2 46.6528
R3 2 N3 30.1089
R4 2 N4 2.3471
R5 2 N5 686.5344m
R6 2 N6 171.2082m
R7 2 N7 40.1594
R8 2 1 10G
R9 2 1 4.1742k
.ends 
*******
.subckt 0402_7447650242_0.42u 1 2
C1 1 N7 19.8327f
L1 1 N1 372.8953n
L2 N1 N2 7.5691n
L3 N2 N3 3.7665n
L4 N3 N4 33.7954n
L5 N4 N5 32.5936n
L6 N5 N6 128.0822n
R1 2 N1 78.5242
R2 2 N2 46.7293
R3 2 N3 30.2765
R4 2 N4 2.3352
R5 2 N5 817.5681m
R6 2 N6 160.0210m
R7 2 N7 40.1594
R8 2 1 10G
R9 2 1 4.5742k
.ends 
*******
.subckt 0402_7447650247_0.47u 1 2
C1 1 N7 24.8327f
L1 1 N1 415.8953n
L2 N1 N2 7.4405n
L3 N2 N3 3.6798n
L4 N3 N4 38.7284n
L5 N4 N5 49.6504n
L6 N5 N6 206.8955n
R1 2 N1 78.4970
R2 2 N2 46.6474
R3 2 N3 30.0979
R4 2 N4 2.3676
R5 2 N5 933.5514m
R6 2 N6 144.8628m
R7 2 N7 40.1594
R8 2 1 10G
R9 2 1 4.4742k
.ends 
*******
.subckt 0402_7447650253_0.53u 1 2
C1 1 N7 16.7711f
L1 1 N1 474n
L2 N1 N2 7.4385n
L3 N2 N3 3.7086n
L4 N3 N4 42.7705n
L5 N4 N5 60.8634n
L6 N5 N6 296.1997n
R1 2 N1 78.4736
R2 2 N2 46.5859
R3 2 N3 29.9610
R4 2 N4 2.3903
R5 2 N5 1.1468
R6 2 N6 112.6878m
R7 2 N7 16.0022
R8 2 1 10g
R9 2 1 5.2773k
.ends 
*******
.subckt 0402_7447650259_0.59u 1 2
C1 1 N7 24.7711f
L1 1 N1 525n
L2 N1 N2 8.4608n
L3 N2 N3 4.7096n
L4 N3 N4 50.1447n
L5 N4 N5 68.0756n
L6 N5 N6 297.6157n
R1 2 N1 78.5427
R2 2 N2 46.8805
R3 2 N3 30.6171
R4 2 N4 2.3824
R5 2 N5 1.3526
R6 2 N6 85.8486m
R7 2 N7 16.0022
R8 2 1 10g
R9 2 1 5.8760k
.ends 
*******
.subckt 0402_7447650270_0.7u 1 2
C1 1 N7 17.7711f
L1 1 N1 635n
L2 N1 N2 7.8439n
L3 N2 N3 4.2048n
L4 N3 N4 53.5064n
L5 N4 N5 146.0545n
L6 N5 N6 637.1949n
R1 2 N1 78.4129
R2 2 N2 46.4883
R3 2 N3 29.7482
R4 2 N4 2.8449
R5 2 N5 1.8006
R6 2 N6 100.8307m
R7 2 N7 16.0022
R8 2 1 10g
R9 2 1 6.2760k
.ends 
*******
.subckt 0402_7447650277_0.77u 1 2
C1 1 N7 25.0598f
L1 1 N1 700n
L2 N1 N2 16.3037n
L3 N2 N3 11.6209n
L4 N3 N4 55.2316n
L5 N4 N5 164.8258n
L6 N5 N6 560.3690n
R1 2 N1 79.3019
R2 2 N2 49.7258
R3 2 N3 36.3877
R4 2 N4 2.9291
R5 2 N5 2.4481
R6 2 N6 16.2631m
R7 2 N7 16.0022
R8 2 1 10g
R9 2 1 8.0760k
.ends 
*******
.subckt 0603_7447610139_0.039u 1 2
C1 1 N7 100.5018f
L1 1 N1 37n
L2 N1 N2 2.0340n
L3 N2 N3 972.6366p
L4 N3 N4 657.9738p
L5 N4 N5 1.5334n
L6 N5 N6 8.1575n
R1 2 N1 239.9382m
R2 2 N2 481.8469m
R3 2 N3 430.1578m
R4 2 N4 314.3276m
R5 2 N5 80.2688m
R6 2 N6 58.6487m
R7 2 N7 3.7517
R8 2 1 10G
R9 2 1 160
.ends 
*******
.subckt 0603_7447610168_0.068u 1 2
C1 1 N7 77.5018f
L1 1 N1 65.8178n
L2 N1 N2 6.4503n
L3 N2 N3 951.1589p
L4 N3 N4 916.7371p
L5 N4 N5 10.7869n
L6 N5 N6 10.0289n
R1 2 N1 394.7042m
R2 2 N2 375.3020m
R3 2 N3 446.7006m
R4 2 N4 365.3678m
R5 2 N5 207.5346m
R6 2 N6 166.1908m
R7 2 N7 100.4162
R8 2 1 10G
R9 2 1 273.7883
.ends 
*******
.subckt 0603_7447610211_0.11u 1 2
C1 1 N7 50.5018f
L1 1 N1 103.8178n
L2 N1 N2 9.2411n
L3 N2 N3 975.8467p
L4 N3 N4 933.6872p
L5 N4 N5 14.7146n
L6 N5 N6 18.7665n
R1 2 N1 867.6254m
R2 2 N2 469.5000m
R3 2 N3 498.3382m
R4 2 N4 416.9726m
R5 2 N5 173.6254m
R6 2 N6 148.4701m
R7 2 N7 100.4162
R8 2 1 10G
R9 2 1 553.7883
.ends 
*******
.subckt 0603_7447610215_0.15u 1 2
C1 1 N7 43.5018f
L1 1 N1 140.8178n
L2 N1 N2 13.2853n
L3 N2 N3 1.0032n
L4 N3 N4 946.4542p
L5 N4 N5 31.1056n
L6 N5 N6 21.9843n
R1 2 N1 1.0309
R2 2 N2 604.9040m
R3 2 N3 566.1729m
R4 2 N4 520.9171m
R5 2 N5 289.3154m
R6 2 N6 303.2085m
R7 2 N7 100.4162
R8 2 1 10G
R9 2 1 689.7883
.ends 
*******
.subckt 0603_7447610220_0.2u 1 2
C1 1 N7 40.5018f
L1 1 N1 211.8178n
L2 N1 N2 17.0122n
L3 N2 N3 9.1407n
L4 N3 N4 1.0475n
L5 N4 N5 54.9967n
L6 N5 N6 65.7191n
R1 2 N1 1.1677
R2 2 N2 668.1253m
R3 2 N3 659.3882m
R4 2 N4 621.7508m
R5 2 N5 390.3418m
R6 2 N6 399.2136m
R7 2 N7 315.0491
R8 2 1 10G
R9 2 1 877.7968
.ends 
*******
.subckt 0603_7447610224_0.24u 1 2
C1 1 N7 58.5018f
L1 1 N1 226.8178n
L2 N1 N2 19.3739n
L3 N2 N3 9.4466n
L4 N3 N4 1.5101n
L5 N4 N5 85.3971n
L6 N5 N6 71.3570n
R1 2 N1 1.9382
R2 2 N2 943.4198m
R3 2 N3 988.0501m
R4 2 N4 975.0542m
R5 2 N5 645.3673m
R6 2 N6 513.2924m
R7 2 N7 15.0491
R8 2 1 10G
R9 2 1 1.2108k
.ends 
*******
.subckt 0603_7447610227_0.27u 1 2
C1 1 N7 39.5018f
L1 1 N1 260n
L2 N1 N2 21.8247n
L3 N2 N3 9.4617n
L4 N3 N4 1.5154n
L5 N4 N5 85.3736n
L6 N5 N6 71.3673n
R1 2 N1 1.9387
R2 2 N2 945.7874m
R3 2 N3 989.1656m
R4 2 N4 976.0803m
R5 2 N5 645.7890m
R6 2 N6 514.1277m
R7 2 N7 15.0491
R8 2 1 10G
R9 2 1 1277.7968
.ends 
*******
.subckt 0603_7447610236_0.36u 1 2
C1 1 N7 65.5018f
L1 1 N1 345n
L2 N1 N2 31.8064n
L3 N2 N3 9.6056n
L4 N3 N4 2.0812n
L5 N4 N5 123.6361n
L6 N5 N6 80.5775n
R1 2 N1 2.7622
R2 2 N2 1.3379
R3 2 N3 1.4017
R4 2 N4 1.3986
R5 2 N5 919.0499m
R6 2 N6 710.5064m
R7 2 N7 15.0491
R8 2 1 10G
R9 2 1 1787.7968
.ends 
*******
.subckt 0603_7447610239_0.39u 1 2
C1 1 N7 70.3088f
L1 1 N1 372n
L2 N1 N2 24.2866n
L3 N2 N3 14.4110n
L4 N3 N4 4.3819n
L5 N4 N5 113.9321n
L6 N5 N6 82.2283n
R1 2 N1 2.8535
R2 2 N2 2.6689
R3 2 N3 2.5266
R4 2 N4 1.2712
R5 2 N5 3097.8744m
R6 2 N6 6360.5101m
R7 2 N7 15.0661
R8 2 1 10G
R9 2 1 1.9630k
.ends 
*******
.subckt 0603_7447610242_0.42u 1 2
C1 1 N7 49.3088f
L1 1 N1 384n
L2 N1 N2 6.4729n
L3 N2 N3 2.8525n
L4 N3 N4 7.0401n
L5 N4 N5 35.4819n
L6 N5 N6 129.9026n
R1 2 N1 78.5206
R2 2 N2 46.6863
R3 2 N3 30.2343
R4 2 N4 2.6817
R5 2 N5 606.0216m
R6 2 N6 669.7126m
R7 2 N7 40.1594
R8 2 1 10G
R9 2 1 1.9630k
.ends 
*******
.subckt 0603_7447610247_0.47u 1 2
C1 1 N7 55.3088f
L1 1 N1 434n
L2 N1 N2 6.1725n
L3 N2 N3 3.0744n
L4 N3 N4 8.0052n
L5 N4 N5 41.8871n
L6 N5 N6 164.3411n
R1 2 N1 78.5121
R2 2 N2 46.7279
R3 2 N3 30.4138
R4 2 N4 3.3308
R5 2 N5 729.4350m
R6 2 N6 466.2101m
R7 2 N7 40.1594
R8 2 1 10G
R9 2 1 2.2130k
.ends 
*******
.subckt 0603_7447610256_0.56u 1 2
C1 1 N7 59.3088f
L1 1 N1 523n
L2 N1 N2 1.2360n
L3 N2 N3 1.5143n
L4 N3 N4 12.5405n
L5 N4 N5 47.1461n
L6 N5 N6 148.0143n
R1 2 N1 78.3268
R2 2 N2 46.4399
R3 2 N3 30.7950
R4 2 N4 4.6396
R5 2 N5 815.7922m
R6 2 N6 604.3792m
R7 2 N7 40.1594
R8 2 1 10G
R9 2 1 2.8930k
.ends 
*******
.subckt 0603_7447610260_0.6u 1 2
C1 1 N7 45.3088f
L1 1 N1 560n
L2 N1 N2 1.0586n
L3 N2 N3 1.3931n
L4 N3 N4 12.7393n
L5 N4 N5 50.8728n
L6 N5 N6 184.1877n
R1 2 N1 78.3255
R2 2 N2 46.4368
R3 2 N3 30.7931
R4 2 N4 4.6564
R5 2 N5 993.7344m
R6 2 N6 604.3792m
R7 2 N7 40.1594
R8 2 1 10G
R9 2 1 2.8330k
.ends 
*******
.subckt 0603_7447610268_0.68u 1 2
C1 1 N7 70.3088f
L1 1 N1 640n
L2 N1 N2 1.0114n
L3 N2 N3 1.3725n
L4 N3 N4 16.0456n
L5 N4 N5 55.6619n
L6 N5 N6 238.0515n
R1 2 N1 78.3246
R2 2 N2 46.4345
R3 2 N3 30.7903
R4 2 N4 4.6674
R5 2 N5 1.0330
R6 2 N6 603.1803m
R7 2 N7 40.1594
R8 2 1 10G
R9 2 1 3.2130k
.ends 
*******
.subckt 0603_7447610282_0.82u 1 2
C1 1 N7 46.3088f
L1 1 N1 775n
L2 N1 N2 983.3826p
L3 N2 N3 1.3957n
L4 N3 N4 26.3384n
L5 N4 N5 68.9543n
L6 N5 N6 307.4580n
R1 2 N1 78.3237
R2 2 N2 46.4326
R3 2 N3 30.7897
R4 2 N4 4.6824
R5 2 N5 1.1502
R6 2 N6 594.8769m
R7 2 N7 300.1594
R8 2 1 10G
R9 2 1 3.8130k
.ends 
*******

.subckt 0603_7447610310_1u 1 2
C1 1 N7 54.3088f
L1 1 N1 945n
L2 N1 N2 981.2366p
L3 N2 N3 1.2999n
L4 N3 N4 44.4258n
L5 N4 N5 88.6737n
L6 N5 N6 577.4982n
R1 2 N1 78.2815
R2 2 N2 46.3122
R3 2 N3 30.5271
R4 2 N4 4.6984
R5 2 N5 1.8128
R6 2 N6 539.3283m
R7 2 N7 300.1594
R8 2 1 10G
R9 2 1 4.9130k
.ends 
*******
.subckt 0603_7447610315_1.5u 1 2
C1 1 N7 46.3088f
L1 1 N1 1.4300u
L2 N1 N2 978.6450p
L3 N2 N3 1.3664n
L4 N3 N4 98.5460n
L5 N4 N5 194.1102n
L6 N5 N6 749.6552n
R1 2 N1 77.9478
R2 2 N2 45.3380
R3 2 N3 28.2081
R4 2 N4 4.7702
R5 2 N5 2.7857
R6 2 N6 432.2827m
R7 2 N7 300.1594
R8 2 1 10G
R9 2 1 7.3130k
.ends 
*******
.subckt 0603_7447610322_2.2u 1 2
C1 1 N7 951.5331f
L1 1 N1 2.1313u
L2 N1 N2 986.1472p
L3 N2 N3 2.2134n
L4 N3 N4 237.1306n
L5 N4 N5 28.2327n
L6 N5 N6 211.4659n
R1 2 N1 77.9937
R2 2 N2 45.4808
R3 2 N3 28.5941
R4 2 N4 4.8281
R5 2 N5 2.2758
R6 2 N6 534.4797m
R7 2 N7 22.4264
R8 2 1 10G
R9 2 1 6.6665k
.ends 
*******
.subckt 0603_7447610333_3.3u 1 2
C1 1 N7 653.3088f
L1 1 N1 3.1900u
L2 N1 N2 987.7903p
L3 N2 N3 2.9628n
L4 N3 N4 290.3709n
L5 N4 N5 670.2000n
L6 N5 N6 1.7729u
R1 2 N1 77.6863
R2 2 N2 44.6101
R3 2 N3 26.7398
R4 2 N4 3.6440
R5 2 N5 3.1695
R6 2 N6 1.1463
R7 2 N7 50.1594
R8 2 1 10G
R9 2 1 10k
.ends 
*******
.subckt 0603_7447610347_4.7u 1 2
C1 1 N7 1.2488p
L1 1 N1 4.5380u
L2 N1 N2 987.0455p
L3 N2 N3 2.9089n
L4 N3 N4 434.8884n
L5 N4 N5 1.4172u
L6 N5 N6 6.4123u
R1 2 N1 77.6177
R2 2 N2 44.3985
R3 2 N3 26.1367
R4 2 N4 4.0412
R5 2 N5 3.2440
R6 2 N6 1.3040
R7 2 N7 2.1594
R8 2 1 10G
R9 2 1 11.3000k
.ends 
*******
.subckt 0603_7447610356_5.6u 1 2
C1 1 N7 1.1988p
L1 1 N1 5.4200u
L2 N1 N2 986.8310p
L3 N2 N3 2.8833n
L4 N3 N4 549.8004n
L5 N4 N5 1.7110u
L6 N5 N6 7.1706u
R1 2 N1 77.5569
R2 2 N2 44.2088
R3 2 N3 25.5719
R4 2 N4 4.1644
R5 2 N5 3.2420
R6 2 N6 1.3800
R7 2 N7 2.1594
R8 2 1 10G
R9 2 1 11.8100k
.ends 
*******
.subckt 0603_7447610368_6.8u 1 2
C1 1 N7 1.4788p
L1 1 N1 6.5600u
L2 N1 N2 986.6500p
L3 N2 N3 2.9572n
L4 N3 N4 708.6023n
L5 N4 N5 2.1614u
L6 N5 N6 14.8928u
R1 2 N1 77.9214
R2 2 N2 45.2740
R3 2 N3 28.4291
R4 2 N4 5.2893
R5 2 N5 3.2941
R6 2 N6 2.0873
R7 2 N7 2.1594
R8 2 1 10G
R9 2 1 13k
.ends 
*******
.subckt 0603_7447610382_8.2u 1 2
C1 1 N7 1.5088p
L1 1 N1 7.8900u
L2 N1 N2 979.4885p
L3 N2 N3 3.2311n
L4 N3 N4 839.2124n
L5 N4 N5 2.7355u
L6 N5 N6 70.2559u
R1 2 N1 80.3420
R2 2 N2 51.8624
R3 2 N3 41.7406
R4 2 N4 5.7739
R5 2 N5 2.9477
R6 2 N6 2.1532
R7 2 N7 2.1577
R8 2 1 10G
R9 2 1 14.4000k
.ends 
*******
.subckt 0603_7447610410_10u 1 2
C1 1 N7 1.7488p
L1 1 N1 9.4900u
L2 N1 N2 977.9088p
L3 N2 N3 3.1164n
L4 N3 N4 1.0174u
L5 N4 N5 3.1179u
L6 N5 N6 99.6612u
R1 2 N1 79.7676
R2 2 N2 50.3739
R3 2 N3 39.3033
R4 2 N4 7.1228
R5 2 N5 2.9437
R6 2 N6 2.1625
R7 2 N7 2.1577
R8 2 1 10G
R9 2 1 15.6200k
.ends 
*******
.subckt 0603_7447610415_15u 1 2
C1 1 N7 1.9788p
L1 1 N1 13.9000u
L2 N1 N2 1.9370n
L3 N2 N3 520.2390n
L4 N3 N4 1.3144u
L5 N4 N5 5.3018u
L6 N5 N6 50.6317u
R1 2 N1 138.6484
R2 2 N2 58.0664
R3 2 N3 67.0319
R4 2 N4 6.7232
R5 2 N5 1.1466
R6 2 N6 1.2249
R7 2 N7 2.1577
R8 2 1 10G
R9 2 1 22.9000k
.ends 
*******
.subckt 0603_7447610422_22u 1 2
C1 1 N7 2.3988p
L1 1 N1 19.1010u
L2 N1 N2 709.8065p
L3 N2 N3 299.9125p
L4 N3 N4 2.2662u
L5 N4 N5 4.8014u
L6 N5 N6 1.4924u
R1 2 N1 106.2913
R2 2 N2 98.9292
R3 2 N3 98.8357
R4 2 N4 8.2048
R5 2 N5 3.0889
R6 2 N6 1.9587
R7 2 N7 2.1124
R8 2 1 10G
R9 2 1 29k
.ends 
*******
.subckt 0805A_744760247A_0.47u 1 2
C1 1 N7 159.5136f
L1 1 N1 450n
L2 N1 N2 20.2094n
L3 N2 N3 18.6247n
L4 N3 N4 583.9523p
L5 N4 N5 9.5844n
L6 N5 N6 1.0575
R1 2 N1 6.1204
R2 2 N2 1.0575
R3 2 N3 9.4334
R4 2 N4 287.0525m
R5 2 N5 8.8470
R6 2 N6 7.1327
R7 2 N7 647.9627
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760256A_0.56u 1 2
C1 1 N7 153.5612f
L1 1 N1 530n
L2 N1 N2 26.8088n
L3 N2 N3 20.2434n
L4 N3 N4 584.2412p
L5 N4 N5 9.5854n
L6 N5 N6 2.4030n
R1 2 N1 6.1191
R2 2 N2 1.0634
R3 2 N3 9.4334
R4 2 N4 294.2585m
R5 2 N5 8.8470
R6 2 N6 7.1327
R7 2 N7 647.5479
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760268A_0.68u 1 2
C1 1 N7 136.6774f
L1 1 N1 663.5n
L2 N1 N2 42.4299n
L3 N2 N3 7.5466n
L4 N3 N4 413.2899p
L5 N4 N5 98.1445n
L6 N5 N6 2.5968n
R1 2 N1 9.4018
R2 2 N2 3.2364
R3 2 N3 9.5397
R4 2 N4 3.3780
R5 2 N5 7.2689
R6 2 N6 8.0843
R7 2 N7 841.5979
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760282A_0.82u 1 2
C1 1 N7 138.9514f
L1 1 N1 770n
L2 N1 N2 8.1508n
L3 N2 N3 2.5651n
L4 N3 N4 40.7889n
L5 N4 N5 14.0322n
L6 N5 N6 12.2484n
R1 2 N1 35.1686
R2 2 N2 18.4937
R3 2 N3 21.2775
R4 2 N4 1.3639
R5 2 N5 9.4796
R6 2 N6 8.0236
R7 2 N7 644.7885
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760310A_1u 1 2
C1 1 N7 127.1422f
L1 1 N1 950n
L2 N1 N2 26.8186n
L3 N2 N3 2.9875n
L4 N3 N4 49.6184n
L5 N4 N5 32.3062n
L6 N5 N6 22.7513n
R1 2 N1 35.2122
R2 2 N2 18.5686
R3 2 N3 21.3253
R4 2 N4 2.5096
R5 2 N5 9.4651
R6 2 N6 7.9994
R7 2 N7 642.5452
R8 2 1 10g
.ends
*******
.subckt 0805A_744760312A_1.2u 1 2
C1 1 N7 127.5473f
L1 1 N1 1.15u
L2 N1 N2 33.5362n
L3 N2 N3 2.6037n
L4 N3 N4 41.1788n
L5 N4 N5 61.5148n
L6 N5 N6 29.7561n
R1 2 N1 37.1888
R2 2 N2 17.7304
R3 2 N3 20.6893
R4 2 N4 2.6032
R5 2 N5 9.4682
R6 2 N6 7.9975
R7 2 N7 697.2085
R8 2 1 10g
.ends 
******* 
.subckt 0805A_744760315A_1.5u 1 2
C1 1 N7 123.1843f
L1 1 N1 1.3757u
L2 N1 N2 57.6285n
L3 N2 N3 3.5418n
L4 N3 N4 55.0942n
L5 N4 N5 49.7480n
L6 N5 N6 31.5411n
R1 2 N1 33.7177
R2 2 N2 20.6069
R3 2 N3 22.8943
R4 2 N4 6.4423
R5 2 N5 9.4804
R6 2 N6 8.0146
R7 2 N7 553.8673
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760318A_1.8u 1 2
C1 1 N7 133.8760f
L1 1 N1 1.65u
L2 N1 N2 65.6086n
L3 N2 N3 3.1064n
L4 N3 N4 60.6754n
L5 N4 N5 79.8796n
L6 N5 N6 40.7869n
R1 2 N1 36.1006
R2 2 N2 21.3755
R3 2 N3 23.5436
R4 2 N4 13.1875
R5 2 N5 9.5493
R6 2 N6 8.1022
R7 2 N7 423.1638
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760322A_2.2u 1 2
C1 1 N7 189.8719f
L1 1 N1 1.8u
L2 N1 N2 450.0742n
L3 N2 N3 2.5035n
L4 N3 N4 5.9638n
L5 N4 N5 7.9713n
L6 N5 N6 4.0616n
R1 2 N1 190.9297
R2 2 N2 24.7252
R3 2 N3 25.7638
R4 2 N4 9.0673
R5 2 N5 9.5964
R6 2 N6 8.1937
R7 2 N7 923.0878
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760327A_2.7u 1 2
C1 1 N7 135.9031f
L1 1 N1 2.25u
L2 N1 N2 583.7325n
L3 N2 N3 3.1043n
L4 N3 N4 6.3162n
L5 N4 N5 8.1769n
L6 N5 N6 4.3153n
R1 2 N1 171.6405
R2 2 N2 24.4242
R3 2 N3 25.4783
R4 2 N4 9.0386
R5 2 N5 9.5704
R6 2 N6 8.1571
R7 2 N7 1.4363k
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760333A_3.3u 1 2
C1 1 N7 158.0233f
L1 1 N1 2.8u
L2 N1 N2 619.9642n
L3 N2 N3 750.4517p
L4 N3 N4 14.5699n
L5 N4 N5 68.6521n
L6 N5 N6 92.0413n
R1 2 N1 157.8926
R2 2 N2 25.8066
R3 2 N3 26.3545
R4 2 N4 26.6522
R5 2 N5 9.8403
R6 2 N6 8.5333
R7 2 N7 1.1054k
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760339A_3.9u 1 2
C1 1 N7 131.1918f
L1 1 N1 3.06u
L2 N1 N2 742.8370n
L3 N2 N3 819.2923p
L4 N3 N4 24.9908n
L5 N4 N5 84.3429n
L6 N5 N6 113.5388n
R1 2 N1 278.1925
R2 2 N2 26.9730
R3 2 N3 27.4690
R4 2 N4 27.9523
R5 2 N5 9.9662
R6 2 N6 8.6837
R7 2 N7 1.3709k
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760347A_4.7u 1 2
C1 1 N7 433.0876f
L1 1 N1 3.9977u
L2 N1 N2 734.0050n
L3 N2 N3 135.2855n
L4 N3 N4 72.2377n
L5 N4 N5 57.2282n
L6 N5 N6 287.7952n
R1 2 N1 198.1838
R2 2 N2 26.0714
R3 2 N3 26.9452
R4 2 N4 27.5069
R5 2 N5 9.8817
R6 2 N6 8.5409
R7 2 N7 784.6283
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760356A_5.6u 1 2
C1 1 N7 459.0344f
L1 1 N1 4.83u
L2 N1 N2 1.0405u
L3 N2 N3 816.1320p
L4 N3 N4 26.4147n
L5 N4 N5 13.1237n
L6 N5 N6 603.8984n
R1 2 N1 218.7445
R2 2 N2 25.3456
R3 2 N3 25.8975
R4 2 N4 26.2602
R5 2 N5 9.7824
R6 2 N6 8.5991
R7 2 N7 486.1824
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760382A_8.2u 1 2
C1 1 N7 291.6740f
L1 1 N1 7.3u
L2 N1 N2 1.2104u
L3 N2 N3 837.1269p
L4 N3 N4 91.4973n
L5 N4 N5 409.6341n
L6 N5 N6 1.3553u
R1 2 N1 272.5206
R2 2 N2 74.3932
R3 2 N3 54.3954
R4 2 N4 56.9118
R5 2 N5 16.4781
R6 2 N6 8.4993
R7 2 N7 851.0096
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760410A_10u 1 2
C1 1 N7 204.4834f
L1 1 N1 8.9u
L2 N1 N2 1.7161u
L3 N2 N3 834.6607p
L4 N3 N4 77.5391n
L5 N4 N5 35.6154n
L6 N5 N6 9.7387u
R1 2 N1 481.9151
R2 2 N2 53.8234
R3 2 N3 53.8243
R4 2 N4 56.4302
R5 2 N5 10.9523
R6 2 N6 8.5315
R7 2 N7 1.1459k
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762312A_1.2u 1 2
C1 1 N7 158.7443f
L1 1 N1 1.15u
L2 N1 N2 25.7595n
L3 N2 N3 2.2471n
L4 N3 N4 35.0721n
L5 N4 N5 49.3056n
L6 N5 N6 26.2082n
R1 2 N1 37.0111
R2 2 N2 16.9448
R3 2 N3 20.1815
R4 2 N4 2.4163
R5 2 N5 9.4612
R6 2 N6 7.9902
R7 2 N7 171.5402
R8 2 1 10g
.ends 
******* 
.subckt 1008A_744762315A_1.5u 1 2
C1 1 N7 144.4482f
L1 1 N1 1.4750u
L2 N1 N2 43.4654n
L3 N2 N3 2.0276n
L4 N3 N4 43.3750n
L5 N4 N5 114.5311n
L6 N5 N6 51.8453n
R1 2 N1 39.7071
R2 2 N2 13.7898
R3 2 N3 18.0981
R4 2 N4 3.2315
R5 2 N5 9.4896
R6 2 N6 8.0124
R7 2 N7 138.0520
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762318A_1.8u 1 2
C1 1 N7 145.4549f
L1 1 N1 1.7850u
L2 N1 N2 57.9562n
L3 N2 N3 3.1587n
L4 N3 N4 9.8599n
L5 N4 N5 68.5705n
L6 N5 N6 27.6903n
R1 2 N1 34.3122
R2 2 N2 20.7754
R3 2 N3 23.0005
R4 2 N4 10.5653
R5 2 N5 9.5416
R6 2 N6 8.1049
R7 2 N7 109.6525
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762322A_2.2u 1 2
C1 1 N7 154.4785f
L1 1 N1 2.16u
L2 N1 N2 76.7015n
L3 N2 N3 4.5985n
L4 N3 N4 11.3131n
L5 N4 N5 72.6643n
L6 N5 N6 26.3276n
R1 2 N1 30.5560
R2 2 N2 21.9301
R3 2 N3 24.0282
R4 2 N4 15.3476
R5 2 N5 9.5424
R6 2 N6 8.1070
R7 2 N7 308.3232
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762327A_2.7u 1 2
C1 1 N7 377.6344f
L1 1 N1 2.65u
L2 N1 N2 120.7859n
L3 N2 N3 3.7238n
L4 N3 N4 7.2030n
L5 N4 N5 9.1192n
L6 N5 N6 4.6590n
R1 2 N1 24.5300
R2 2 N2 23.4744
R3 2 N3 29.1481
R4 2 N4 29.7704
R5 2 N5 20.5211
R6 2 N6 8.5261
R7 2 N7 172.7902
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762333A_3.3u 1 2
C1 1 N7 511.8368f
L1 1 N1 3.1u
L2 N1 N2 301.2330n
L3 N2 N3 744.1133p
L4 N3 N4 38.9127n
L5 N4 N5 47.9265n
L6 N5 N6 204.2512n
R1 2 N1 277.7959
R2 2 N2 26.2115
R3 2 N3 26.7451
R4 2 N4 27.1918
R5 2 N5 9.8920
R6 2 N6 8.5597
R7 2 N7 56.1459
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762339A_3.9u 1 2
C1 1 N7 713.2456f
L1 1 N1 3.6u
L2 N1 N2 182.3549n
L3 N2 N3 757.0463p
L4 N3 N4 139.0604n
L5 N4 N5 45.5489n
L6 N5 N6 2.0109u
R1 2 N1 142.0736
R2 2 N2 28.2253
R3 2 N3 28.6967
R4 2 N4 20.2129
R5 2 N5 9.9985
R6 2 N6 18.6399
R7 2 N7 135.2796
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762347A_4.7u 1 2
C1 1 N7 702.5978f
L1 1 N1 4.45u
L2 N1 N2 248.4266n
L3 N2 N3 757.2336p
L4 N3 N4 127.8327n
L5 N4 N5 51.0308n
L6 N5 N6 651.0043n
R1 2 N1 159.2400
R2 2 N2 28.7319
R3 2 N3 26.2849
R4 2 N4 25.4177
R5 2 N5 16.2226
R6 2 N6 19.2937
R7 2 N7 156.4933
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762356A_5.6u 1 2
C1 1 N7 323.8953f
L1 1 N1 5.1u
L2 N1 N2 605.4820n
L3 N2 N3 757.3560p
L4 N3 N4 327.1355n
L5 N4 N5 50.1316n
L6 N5 N6 588.7510n
R1 2 N1 185.5893
R2 2 N2 28.7002
R3 2 N3 26.2381
R4 2 N4 26.1783
R5 2 N5 18.6959
R6 2 N6 20.8881
R7 2 N7 268.1882
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762368A_6.8u 1 2
C1 1 N7 500.1575f
L1 1 N1 6.1u
L2 N1 N2 860.1723n
L3 N2 N3 761.1966p
L4 N3 N4 56.2783n
L5 N4 N5 59.2882n
L6 N5 N6 1.1711u
R1 2 N1 262.2656
R2 2 N2 30.7085
R3 2 N3 28.5802
R4 2 N4 28.9585
R5 2 N5 23.5813
R6 2 N6 21.3351
R7 2 N7 146.3916
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762382A_8.2u 1 2
C1 1 N7 730.0597f
L1 1 N1 7.25u
L2 N1 N2 962.4842n
L3 N2 N3 762.2250p
L4 N3 N4 60.3358n
L5 N4 N5 61.7402n
L6 N5 N6 2.2536u
R1 2 N1 265.8819
R2 2 N2 31.4736
R3 2 N3 29.4515
R4 2 N4 29.7693
R5 2 N5 24.4361
R6 2 N6 21.2667
R7 2 N7 127.7118
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762410A_10u 1 2
C1 1 N7 855.8897f
L1 1 N1 8.9u
L2 N1 N2 1.1434u
L3 N2 N3 762.6593p
L4 N3 N4 62.6732n
L5 N4 N5 63.2942n
L6 N5 N6 2.9201u
R1 2 N1 270.7618
R2 2 N2 32.1396
R3 2 N3 30.2058
R4 2 N4 30.4913
R5 2 N5 25.4603
R6 2 N6 21.1285
R7 2 N7 145.5541
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762415A_15u 1 2
C1 1 N7 365.0719f
L1 1 N1 14u
L2 N1 N2 2.6334u
L3 N2 N3 834.7144p
L4 N3 N4 77.5391n
L5 N4 N5 36.3963n
L6 N5 N6 9.8862u
R1 2 N1 558.8531
R2 2 N2 74.1014
R3 2 N3 64.1023
R4 2 N4 76.6831
R5 2 N5 21.3423
R6 2 N6 48.5308
R7 2 N7 109.0096
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762418A_18u 1 2
C1 1 N7 1.7966p
L1 1 N1 16.9u
L2 N1 N2 1.2439u
L3 N2 N3 836.0875p
L4 N3 N4 837.1967p
L5 N4 N5 269.6004n
L6 N5 N6 9.6504u
R1 2 N1 88.8571
R2 2 N2 55.2375
R3 2 N3 55.2405
R4 2 N4 25.7197
R5 2 N5 49.3684
R6 2 N6 18.5307
R7 2 N7 199.5243
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762422A_22u 1 2
C1 1 N7 564.1908f
L1 1 N1 20u
L2 N1 N2 2.2755u
L3 N2 N3 834.6409p
L4 N3 N4 834.7236p
L5 N4 N5 42.0581n
L6 N5 N6 1.2318u
R1 2 N1 339.4305
R2 2 N2 135.6962
R3 2 N3 133.7892
R4 2 N4 91.0732
R5 2 N5 36.1596
R6 2 N6 77.1113
R7 2 N7 264.3824
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762427A_27u 1 2
C1 1 N7 842.5091f
L1 1 N1 25u
L2 N1 N2 2.5507u
L3 N2 N3 835.3527p
L4 N3 N4 835.4006p
L5 N4 N5 42.3375n
L6 N5 N6 7.3808u
R1 2 N1 374.3260
R2 2 N2 259.8700
R3 2 N3 158.2613
R4 2 N4 130.9240
R5 2 N5 39.7641
R6 2 N6 126.2110
R7 2 N7 249.3839
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762433A_33u 1 2
C1 1 N7 887.1570f
L1 1 N1 30.3u
L2 N1 N2 3.1301u
L3 N2 N3 836.3149p
L4 N3 N4 836.3629p
L5 N4 N5 42.7424n
L6 N5 N6 7.6794u
R1 2 N1 371.5537
R2 2 N2 260.7929
R3 2 N3 160.6972
R4 2 N4 134.4474
R5 2 N5 40.1332
R6 2 N6 125.9908
R7 2 N7 228.6092
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762439A_39u 1 2
C1 1 N7 749.6654f
L1 1 N1 34.7u
L2 N1 N2 4.6998u
L3 N2 N3 835.9555p
L4 N3 N4 836.0075p
L5 N4 N5 43.6164n
L6 N5 N6 9.7186u
R1 2 N1 358.9162
R2 2 N2 267.3951
R3 2 N3 267.4135
R4 2 N4 177.2095
R5 2 N5 45.8166
R6 2 N6 127.5346
R7 2 N7 209.5201
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762447A_47u 1 2
C1 1 N7 619.3667f
L1 1 N1 43.7u
L2 N1 N2 3.3960u
L3 N2 N3 836.2281p
L4 N3 N4 836.3151p
L5 N4 N5 46.4124n
L6 N5 N6 32.0350u
R1 2 N1 341.5274
R2 2 N2 294.2093
R3 2 N3 294.2254
R4 2 N4 235.2256
R5 2 N5 54.7054
R6 2 N6 129.2261
R7 2 N7 292.1897
R8 2 1 10g
.ends 
*******