**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Power Inductor
* Matchcode:              WE-PD4
* Library Type:           spice
* Version:                rev
* Created/modified by:    Ella
* Date and Time:          7/12/2024
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
.subckt TypeL_7445601_1u 1 2
Rp 1 2 2750
Cp 1 2 3.5p
Rs 1 N3 0.004
L1 N3 2 0.803u
.ends TypeL_7445601_1u
*******
.subckt TypeL_74456015_1.5u 1 2
Rp 1 2 4200
Cp 1 2 4p
Rs 1 N3 0.006
L1 N3 2 1.1u
.ends TypeL_74456015_1.5u
*******
.subckt TypeL_74456022_2.2u 1 2
Rp 1 2 7100
Cp 1 2 3p
Rs 1 N3 0.007
L1 N3 2 1.95u
.ends TypeL_74456022_2.2u
*******
.subckt TypeL_74456025_2.5u 1 2
Rp 1 2 7100
Cp 1 2 4.8p
Rs 1 N3 0.009
L1 N3 2 2u
.ends TypeL_74456025_2.5u
*******
.subckt TypeL_74456033_3.3u 1 2
Rp 1 2 7700
Cp 1 2 5.2p
Rs 1 N3 0.011
L1 N3 2 2.6u
.ends TypeL_74456033_3.3u
*******
.subckt TypeL_74456047_4.7u 1 2
Rp 1 2 10150
Cp 1 2 5.2p
Rs 1 N3 0.015
L1 N3 2 3.7u
.ends TypeL_74456047_4.7u
*******
.subckt TypeL_74456056_5.6u 1 2
Rp 1 2 12850
Cp 1 2 6p
Rs 1 N3 0.024
L1 N3 2 4.8u
.ends TypeL_74456056_5.6u
*******
.subckt TypeL_74456068_6.8u 1 2
Rp 1 2 15200
Cp 1 2 4.75p
Rs 1 N3 0.026
L1 N3 2 5.8u
.ends TypeL_74456068_6.8u
*******
.subckt TypeL_74456082_8.2u 1 2
Rp 1 2 15500
Cp 1 2 5.5p
Rs 1 N3 0.034
L1 N3 2 6.8u
.ends TypeL_74456082_8.2u
*******
.subckt TypeL_7445610_10u 1 2
Rp 1 2 18300
Cp 1 2 5.5p
Rs 1 N3 0.035
L1 N3 2 8.35u
.ends TypeL_7445610_10u
*******
.subckt TypeL_74456115_15u 1 2
Rp 1 2 23920
Cp 1 2 6.6p
Rs 1 N3 0.043
L1 N3 2 12.9u
.ends TypeL_74456115_15u
*******
.subckt TypeL_74456122_22u 1 2
Rp 1 2 34700
Cp 1 2 6.25p
Rs 1 N3 0.071
L1 N3 2 19.1u
.ends TypeL_74456122_22u
*******
.subckt TypeL_74456133_33u 1 2
Rp 1 2 40000
Cp 1 2 5.8p
Rs 1 N3 0.094
L1 N3 2 26.5u
.ends TypeL_74456133_33u
*******
.subckt TypeL_74456147_47u 1 2
Rp 1 2 55600
Cp 1 2 5.9p
Rs 1 N3 0.142
L1 N3 2 39.15u
.ends TypeL_74456147_47u
*******
.subckt TypeL_74456168_68u 1 2
Rp 1 2 58200
Cp 1 2 5.4p
Rs 1 N3 0.187
L1 N3 2 58.2u
.ends TypeL_74456168_68u
*******
.subckt TypeL_7445620_100u 1 2
Rp 1 2 80000
Cp 1 2 6.6p
Rs 1 N3 0.253
L1 N3 2 82.35u
.ends TypeL_7445620_100u
*******
.subckt TypeL_74456215_150u 1 2
Rp 1 2 89500
Cp 1 2 6.7p
Rs 1 N3 0.448
L1 N3 2 129.5u
.ends TypeL_74456215_150u
*******
.subckt TypeL_74456222_220u 1 2
Rp 1 2 94000
Cp 1 2 6p
Rs 1 N3 0.601
L1 N3 2 187.5u
.ends TypeL_74456222_220u
*******
.subckt TypeL_74456233_330u 1 2
Rp 1 2 94700
Cp 1 2 6p
Rs 1 N3 0.893
L1 N3 2 276.75u
.ends TypeL_74456233_330u
*******
.subckt TypeL_74456247_470u 1 2
Rp 1 2 125100
Cp 1 2 6.3p
Rs 1 N3 1.315
L1 N3 2 412.15u
.ends TypeL_74456247_470u
*******
.subckt TypeL_74456268_680u 1 2
Rp 1 2 140950
Cp 1 2 7.7p
Rs 1 N3 1.942
L1 N3 2 600u
.ends TypeL_74456268_680u
*******
.subckt TypeL_7445630_1000u 1 2
Rp 1 2 160500
Cp 1 2 8.1p
Rs 1 N3 2.94
L1 N3 2 901u
.ends TypeL_7445630_1000u
*******
.subckt TypeL_74456322_2200u 1 2
Rp 1 2 235150
Cp 1 2 8.9p
Rs 1 N3 6.26
L1 N3 2 1800u
.ends TypeL_74456322_2200u
*******
.subckt TypeL_74456347_4700u 1 2
Rp 1 2 278200
Cp 1 2 6.94p
Rs 1 N3 13.3
L1 N3 2 4200u
.ends TypeL_74456347_4700u
*******
.subckt TypeL_74456382_8200u 1 2
Rp 1 2 848000
Cp 1 2 7.4p
Rs 1 N3 28
L1 N3 2 6250u
.ends TypeL_74456382_8200u
*******
.subckt TypeL_7445640_10000u 1 2
Rp 1 2 1620000
Cp 1 2 6.7p
Rs 1 N3 29.9
L1 N3 2 9000u
.ends TypeL_7445640_10000u
*******
.subckt TypeS_7445501_1u 1 2
Rp 1 2 1100
Cp 1 2 5.9p
Rs 1 N3 0.017
L1 N3 2 0.8u
.ends TypeS_7445501_1u
*******
.subckt TypeS_74455015_1.5u 1 2
Rp 1 2 2350
Cp 1 2 4.5p
Rs 1 N3 0.02
L1 N3 2 1.3u
.ends TypeS_74455015_1.5u
*******
.subckt TypeS_74455022_2.2u 1 2
Rp 1 2 2650
Cp 1 2 3.85p
Rs 1 N3 0.028
L1 N3 2 2.2u
.ends TypeS_74455022_2.2u
*******
.subckt TypeS_74455033_3.3u 1 2
Rp 1 2 2800
Cp 1 2 5.5p
Rs 1 N3 0.044
L1 N3 2 3u
.ends TypeS_74455033_3.3u
*******
.subckt TypeS_74455047_4.7u 1 2
Rp 1 2 5600
Cp 1 2 4.7p
Rs 1 N3 0.063
L1 N3 2 3.75u
.ends TypeS_74455047_4.7u
*******
.subckt TypeS_74455068_6.8u 1 2
Rp 1 2 8500
Cp 1 2 5.45p
Rs 1 N3 0.092
L1 N3 2 5.7u
.ends TypeS_74455068_6.8u
*******
.subckt TypeS_7445510_10u 1 2
Rp 1 2 9700
Cp 1 2 4p
Rs 1 N3 0.121
L1 N3 2 9.1u
.ends TypeS_7445510_10u
*******
.subckt TypeS_74455115_15u 1 2
Rp 1 2 13600
Cp 1 2 5.8p
Rs 1 N3 0.176
L1 N3 2 11.7u
.ends TypeS_74455115_15u
*******
.subckt TypeS_74455122_22u 1 2
Rp 1 2 23200
Cp 1 2 5.6p
Rs 1 N3 0.255
L1 N3 2 18.6u
.ends TypeS_74455122_22u
*******
.subckt TypeS_74455133_33u 1 2
Rp 1 2 33000
Cp 1 2 4.8p
Rs 1 N3 0.362
L1 N3 2 27.2u
.ends TypeS_74455133_33u
*******
.subckt TypeS_74455147_47u 1 2
Rp 1 2 33000
Cp 1 2 4.2p
Rs 1 N3 0.556
L1 N3 2 41.6u
.ends TypeS_74455147_47u
*******
.subckt TypeS_74455168_68u 1 2
Rp 1 2 38500
Cp 1 2 5.1p
Rs 1 N3 0.79
L1 N3 2 51.6u
.ends TypeS_74455168_68u
*******
.subckt TypeS_7445520_100u 1 2
Rp 1 2 52800
Cp 1 2 4.5p
Rs 1 N3 1.08
L1 N3 2 86u
.ends TypeS_7445520_100u
*******
.subckt TypeS_74455215_150u 1 2
Rp 1 2 53100
Cp 1 2 5.65p
Rs 1 N3 1.45
L1 N3 2 135u
.ends TypeS_74455215_150u
*******
.subckt TypeS_74455222_220u 1 2
Rp 1 2 79250
Cp 1 2 5.35p
Rs 1 N3 2.58
L1 N3 2 197u
.ends TypeS_74455222_220u
*******
.subckt TypeS_74455233_330u 1 2
Rp 1 2 128600
Cp 1 2 5.4p
Rs 1 N3 4.15
L1 N3 2 292u
.ends TypeS_74455233_330u
*******
.subckt TypeS_74455247_470u 1 2
Rp 1 2 138000
Cp 1 2 6.45p
Rs 1 N3 5.58
L1 N3 2 401.4u
.ends TypeS_74455247_470u
*******
.subckt TypeS_7445530_1000u 1 2
Rp 1 2 253250
Cp 1 2 6p
Rs 1 N3 11.5
L1 N3 2 814.9u
.ends TypeS_7445530_1000u
*******
.subckt TypeX_74458001_1u 1 2
Rp 1 2 798
Cp 1 2 5.4p
Rs 1 N3 0.005
L1 N3 2 0.85u
.ends TypeX_74458001_1u
*******
.subckt TypeX_74458002_2.2u 1 2
Rp 1 2 1100
Cp 1 2 7.2p
Rs 1 N3 0.008
L1 N3 2 2u
.ends TypeX_74458002_2.2u
*******
.subckt TypeX_74458003_3.3u 1 2
Rp 1 2 2780
Cp 1 2 8.2p
Rs 1 N3 0.01
L1 N3 2 2.8u
.ends TypeX_74458003_3.3u
*******
.subckt TypeX_74458005_5.6u 1 2
Rp 1 2 4680
Cp 1 2 8.5p
Rs 1 N3 0.012
L1 N3 2 4.5u
.ends TypeX_74458005_5.6u
*******
.subckt TypeX_74458010_10u 1 2
Rp 1 2 9200
Cp 1 2 6.5p
Rs 1 N3 0.021
L1 N3 2 8.5u
.ends TypeX_74458010_10u
*******
.subckt TypeX_74458115_15u 1 2
Rp 1 2 13700
Cp 1 2 8.5p
Rs 1 N3 0.03
L1 N3 2 12.1u
.ends TypeX_74458115_15u
*******
.subckt TypeX_74458122_22u 1 2
Rp 1 2 18700
Cp 1 2 7.7p
Rs 1 N3 0.043
L1 N3 2 18.5u
.ends TypeX_74458122_22u
*******
.subckt TypeX_74458133_33u 1 2
Rp 1 2 29200
Cp 1 2 8.6p
Rs 1 N3 0.06
L1 N3 2 27.6u
.ends TypeX_74458133_33u
*******
.subckt TypeX_74458147_47u 1 2
Rp 1 2 34500
Cp 1 2 9p
Rs 1 N3 0.076
L1 N3 2 39.15u
.ends TypeX_74458147_47u
*******
.subckt TypeX_74458168_68u 1 2
Rp 1 2 41900
Cp 1 2 9p
Rs 1 N3 0.11
L1 N3 2 58.75u
.ends TypeX_74458168_68u
*******
.subckt TypeX_7445820_100u 1 2
Rp 1 2 57500
Cp 1 2 7.7p
Rs 1 N3 0.141
L1 N3 2 80.1u
.ends TypeX_7445820_100u
*******
.subckt TypeX_74458215_150u 1 2
Rp 1 2 67600
Cp 1 2 9.4p
Rs 1 N3 0.21
L1 N3 2 116.15u
.ends TypeX_74458215_150u
*******
.subckt TypeX_74458220_220u 1 2
Rp 1 2 71000
Cp 1 2 13p
Rs 1 N3 0.326
L1 N3 2 183u
.ends TypeX_74458220_220u
*******
.subckt TypeX_74458233_330u 1 2
Rp 1 2 74400
Cp 1 2 13p
Rs 1 N3 0.431
L1 N3 2 274u
.ends TypeX_74458233_330u
*******
.subckt TypeX_74458247_470u 1 2
Rp 1 2 90300
Cp 1 2 13p
Rs 1 N3 0.633
L1 N3 2 379.6u
.ends TypeX_74458247_470u
*******
.subckt TypeX_74458268_680u 1 2
Rp 1 2 102100
Cp 1 2 13.2p
Rs 1 N3 0.954
L1 N3 2 592.3u
.ends TypeX_74458268_680u
*******
.subckt TypeX_7445830_1000u 1 2
Rp 1 2 103800
Cp 1 2 14.15p
Rs 1 N3 1.37
L1 N3 2 778.3u
.ends TypeX_7445830_1000u
*******
.subckt TypeXL_74457006_0.5u 1 2
Rp 1 2 2100
Cp 1 2 4.6p
Rs 1 N3 0.001
L1 N3 2 0.4u
.ends TypeXL_74457006_0.5u
*******
.subckt TypeXL_74457008_0.8u 1 2
Rp 1 2 2900
Cp 1 2 4.6p
Rs 1 N3 0.002
L1 N3 2 0.41u
.ends TypeXL_74457008_0.8u
*******
.subckt TypeXL_74457010_1u 1 2
Rp 1 2 3900
Cp 1 2 3.7p
Rs 1 N3 0.003
L1 N3 2 0.8u
.ends TypeXL_74457010_1u
*******
.subckt TypeXL_74457012_1.2u 1 2
Rp 1 2 5500
Cp 1 2 4.95p
Rs 1 N3 0.003
L1 N3 2 1.1u
.ends TypeXL_74457012_1.2u
*******
.subckt TypeXL_74457018_1.8u 1 2
Rp 1 2 6400
Cp 1 2 5.1p
Rs 1 N3 0.005
L1 N3 2 1.7u
.ends TypeXL_74457018_1.8u
*******
.subckt TypeXL_74457027_2.7u 1 2
Rp 1 2 7100
Cp 1 2 5.2p
Rs 1 N3 0.007
L1 N3 2 2.5u
.ends TypeXL_74457027_2.7u
*******
.subckt TypeXL_74457033_3.3u 1 2
Rp 1 2 12100
Cp 1 2 5.5p
Rs 1 N3 0.008
L1 N3 2 3u
.ends TypeXL_74457033_3.3u
*******
.subckt TypeXL_74457047_4.7u 1 2
Rp 1 2 13500
Cp 1 2 6.5p
Rs 1 N3 0.009
L1 N3 2 3.7u
.ends TypeXL_74457047_4.7u
*******
.subckt TypeXL_74457056_5.6u 1 2
Rp 1 2 12000
Cp 1 2 6p
Rs 1 N3 0.012
L1 N3 2 4.8u
.ends TypeXL_74457056_5.6u
*******
.subckt TypeXL_74457068_6.8u 1 2
Rp 1 2 17500
Cp 1 2 6.3p
Rs 1 N3 0.014
L1 N3 2 6u
.ends TypeXL_74457068_6.8u
*******
.subckt TypeXL_74457082_8.2u 1 2
Rp 1 2 20400
Cp 1 2 7.1p
Rs 1 N3 0.016
L1 N3 2 6.8u
.ends TypeXL_74457082_8.2u
*******
.subckt TypeXL_7445710_10u 1 2
Rp 1 2 20700
Cp 1 2 6.6p
Rs 1 N3 0.017
L1 N3 2 7.8u
.ends TypeXL_7445710_10u
*******
.subckt TypeXL_74457112_12u 1 2
Rp 1 2 24500
Cp 1 2 6.6p
Rs 1 N3 0.024
L1 N3 2 10u
.ends TypeXL_74457112_12u
*******
.subckt TypeXL_74457115_15u 1 2
Rp 1 2 19200
Cp 1 2 8.1p
Rs 1 N3 0.029
L1 N3 2 12.7u
.ends TypeXL_74457115_15u
*******
.subckt TypeXL_74457118_18u 1 2
Rp 1 2 32500
Cp 1 2 6.7p
Rs 1 N3 0.033
L1 N3 2 15u
.ends TypeXL_74457118_18u
*******
.subckt TypeXL_74457122_22u 1 2
Rp 1 2 35500
Cp 1 2 7.4p
Rs 1 N3 0.039
L1 N3 2 18u
.ends TypeXL_74457122_22u
*******
.subckt TypeXL_74457127_27u 1 2
Rp 1 2 37200
Cp 1 2 7.5p
Rs 1 N3 0.044
L1 N3 2 21.65u
.ends TypeXL_74457127_27u
*******
.subckt TypeXL_74457133_33u 1 2
Rp 1 2 37400
Cp 1 2 7.6p
Rs 1 N3 0.058
L1 N3 2 26.2u
.ends TypeXL_74457133_33u
*******
.subckt TypeXL_74457139_39u 1 2
Rp 1 2 45400
Cp 1 2 7.15p
Rs 1 N3 0.065
L1 N3 2 31.3u
.ends TypeXL_74457139_39u
*******
.subckt TypeXL_74457147_47u 1 2
Rp 1 2 48400
Cp 1 2 8.3p
Rs 1 N3 0.091
L1 N3 2 39.6u
.ends TypeXL_74457147_47u
*******
.subckt TypeXL_74457156_56u 1 2
Rp 1 2 52600
Cp 1 2 7.7p
Rs 1 N3 0.097
L1 N3 2 45.1u
.ends TypeXL_74457156_56u
*******
.subckt TypeXL_74457168_68u 1 2
Rp 1 2 53800
Cp 1 2 7.8p
Rs 1 N3 0.112
L1 N3 2 56.2u
.ends TypeXL_74457168_68u
*******
.subckt TypeXL_74457182_82u 1 2
Rp 1 2 62650
Cp 1 2 7.6p
Rs 1 N3 0.144
L1 N3 2 68.8u
.ends TypeXL_74457182_82u
*******
.subckt TypeXL_7445720_100u 1 2
Rp 1 2 66400
Cp 1 2 7.8p
Rs 1 N3 0.168
L1 N3 2 78.5u
.ends TypeXL_7445720_100u
*******
.subckt TypeXL_74457212_120u 1 2
Rp 1 2 63500
Cp 1 2 12.6p
Rs 1 N3 0.196
L1 N3 2 108.3u
.ends TypeXL_74457212_120u
*******
.subckt TypeXL_74457215_150u 1 2
Rp 1 2 63550
Cp 1 2 11.7p
Rs 1 N3 0.223
L1 N3 2 125.1u
.ends TypeXL_74457215_150u
*******
.subckt TypeXL_74457218_180u 1 2
Rp 1 2 59900
Cp 1 2 12p
Rs 1 N3 0.256
L1 N3 2 153u
.ends TypeXL_74457218_180u
*******
.subckt TypeXL_74457222_220u 1 2
Rp 1 2 61500
Cp 1 2 12.3p
Rs 1 N3 0.323
L1 N3 2 178.9u
.ends TypeXL_74457222_220u
*******
.subckt TypeXL_74457227_270u 1 2
Rp 1 2 73700
Cp 1 2 13p
Rs 1 N3 0.399
L1 N3 2 228u
.ends TypeXL_74457227_270u
*******
.subckt TypeXL_74457230_1000u 1 2
Rp 1 2 95100
Cp 1 2 12.6p
Rs 1 N3 1.506
L1 N3 2 899u
.ends TypeXL_74457230_1000u
*******
.subckt TypeXL_74457233_330u 1 2
Rp 1 2 74100
Cp 1 2 13.7p
Rs 1 N3 0.47
L1 N3 2 278.5u
.ends TypeXL_74457233_330u
*******
.subckt TypeXL_74457239_390u 1 2
Rp 1 2 74300
Cp 1 2 12.2p
Rs 1 N3 0.558
L1 N3 2 326.7u
.ends TypeXL_74457239_390u
*******
.subckt TypeXL_74457247_470u 1 2
Rp 1 2 79700
Cp 1 2 12.5p
Rs 1 N3 0.674
L1 N3 2 417.7u
.ends TypeXL_74457247_470u
*******
.subckt TypeXL_74457256_560u 1 2
Rp 1 2 79400
Cp 1 2 13.6p
Rs 1 N3 0.855
L1 N3 2 476.5u
.ends TypeXL_74457256_560u
*******
.subckt TypeXL_74457268_680u 1 2
Rp 1 2 81500
Cp 1 2 13.2p
Rs 1 N3 1.002
L1 N3 2 548.3u
.ends TypeXL_74457268_680u
*******
.subckt TypeXL_74457282_820u 1 2
Rp 1 2 93200
Cp 1 2 14.2p
Rs 1 N3 1.172
L1 N3 2 622.5u
.ends TypeXL_74457282_820u
*******
