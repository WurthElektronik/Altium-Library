**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Shielded Coupled Inductor
* Matchcode:              WE-DD 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1210_7448709022_2.2u  1  2  3  4  PARAMS:
+  Cww=15.397p
+  Rp1=4571.89909972
+  Cp1=4.377137093905p
+  Lp1=2.04254489984u
+  Rp2=4571.89909972
+  Cp2=4.377137093905p
+  Lp2=2.04254489984u
+  RDC1=1.67500004172325E-02
+  RDC2=1.67500004172325E-02
+  K=0.93166089804381
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1210_7448709033_3.3u  1  2  3  4  PARAMS:
+  Cww=16.758p
+  Rp1=5734.002646107
+  Cp1=4.826841480055p
+  Lp1=2.871069399387u
+  Rp2=5734.002646107
+  Cp2=4.826841480055p
+  Lp2=2.871069399387u
+  RDC1=0.018499999307096
+  RDC2=0.018499999307096
+  K=0.948495190413777
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1210_7448709047_4.7u  1  2  3  4  PARAMS:
+  Cww=17.045p
+  Rp1=7323.889458193
+  Cp1=6.320129473245p
+  Lp1=3.653348053149u
+  Rp2=7323.889458193
+  Cp2=6.320129473245p
+  Lp2=3.653348053149u
+  RDC1=0.019749999511987
+  RDC2=0.019749999511987
+  K=0.924393723985322
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1210_7448709068_6.8u  1  2  3  4  PARAMS:
+  Cww=22.053p
+  Rp1=8686.592099699
+  Cp1=10.370323770498p
+  Lp1=6.044956452362u
+  Rp2=8686.592099699
+  Cp2=10.370323770498p
+  Lp2=6.044956452362u
+  RDC1=2.27500000037253E-02
+  RDC2=2.27500000037253E-02
+  K=0.957483236357168
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1210_7448709100_10u  1  2  3  4  PARAMS:
+  Cww=19.605p
+  Rp1=15108.50684971
+  Cp1=4.809452174944p
+  Lp1=9.092163844674u
+  Rp2=15108.50684971
+  Cp2=4.809452174944p
+  Lp2=9.092163844674u
+  RDC1=3.20000001229346E-02
+  RDC2=3.20000001229346E-02
+  K=0.965028354684641
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1210_7448709220_22u  1  2  3  4  PARAMS:
+  Cww=27.985p
+  Rp1=22274.55537681
+  Cp1=10.192199908148p
+  Lp1=18.67311530234u
+  Rp2=22274.55537681
+  Cp2=10.192199908148p
+  Lp2=18.67311530234u
+  RDC1=6.35000001639128E-02
+  RDC2=6.35000001639128E-02
+  K=0.970093458055336
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1210_7448709330_33u  1  2  3  4  PARAMS:
+  Cww=32.37p
+  Rp1=24284.43136206
+  Cp1=21.00908036781p
+  Lp1=28.81007759381u
+  Rp2=24284.43136206
+  Cp2=21.00908036781p
+  Lp2=28.81007759381u
+  RDC1=8.15000012516975E-02
+  RDC2=8.15000012516975E-02
+  K=0.969081540939246
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1210_7448709470_47u  1  2  3  4  PARAMS:
+  Cww=32.925p
+  Rp1=25379.79072803
+  Cp1=35.25875980975p
+  Lp1=39.47609509549u
+  Rp2=25379.79072803
+  Cp2=35.25875980975p
+  Lp2=39.47609509549u
+  RDC1=0.106000000610948
+  RDC2=0.106000000610948
+  K=0.970071567724498
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744871004_4.7u  1  2  3  4  PARAMS:
+  Cww=8.435p
+  Rp1=6466.134965155
+  Cp1=10.474822618877p
+  Lp1=3.73454586566u
+  Rp2=6466.134965155
+  Cp2=10.474822618877p
+  Lp2=3.73454586566u
+  RDC1=2.17499998398125E-02
+  RDC2=2.17499998398125E-02
+  K=0.923497267759563
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744871006_6.8u  1  2  3  4  PARAMS:
+  Cww=11.86p
+  Rp1=9328.218597861
+  Cp1=13.421191062565p
+  Lp1=5.912058604035u
+  Rp2=9328.218597861
+  Cp2=13.421191062565p
+  Lp2=5.912058604035u
+  RDC1=0.029250000603497
+  RDC2=0.029250000603497
+  K=0.932857144336311
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744871101_100u  1  2  3  4  PARAMS:
+  Cww=19.08p
+  Rp1=68675.31663075
+  Cp1=23.05282500058p
+  Lp1=78.72494041094u
+  Rp2=68675.31663075
+  Cp2=23.05282500058p
+  Lp2=78.72494041094u
+  RDC1=0.254249997437
+  RDC2=0.254249997437
+  K=0.933112129244154
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744871220_22u  1  2  3  4  PARAMS:
+  Cww=11.51p
+  Rp1=22638.73967817
+  Cp1=15.11440936641p
+  Lp1=18.3534998017u
+  Rp2=22638.73967817
+  Cp2=15.11440936641p
+  Lp2=18.3534998017u
+  RDC1=6.65000006556511E-02
+  RDC2=6.65000006556511E-02
+  K=0.916852926963767
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744871330_33u  1  2  3  4  PARAMS:
+  Cww=10.09p
+  Rp1=37975.78013716
+  Cp1=15.75831604781p
+  Lp1=27.42134037793u
+  Rp2=37975.78013716
+  Cp2=15.75831604781p
+  Lp2=27.42134037793u
+  RDC1=0.10050000064075
+  RDC2=0.10050000064075
+  K=0.930766843975673
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744871470_47u  1  2  3  4  PARAMS:
+  Cww=12.6p
+  Rp1=34885.54369855
+  Cp1=22.22568355332p
+  Lp1=38.57634631342u
+  Rp2=34885.54369855
+  Cp2=22.22568355332p
+  Lp2=38.57634631342u
+  RDC1=0.152000002563
+  RDC2=0.152000002563
+  K=0.925190486042731
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874001_1.5u  1  2  3  4  PARAMS:
+  Cww=14.33p
+  Rp1=3588.593577704
+  Cp1=3.43458631932p
+  Lp1=1.480304877396u
+  Rp2=3588.593577704
+  Cp2=3.43458631932p
+  Lp2=1.480304877396u
+  RDC1=1.25750000588596E-02
+  RDC2=1.25750000588596E-02
+  K=0.967824967992805
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874002_2.4u  1  2  3  4  PARAMS:
+  Cww=12.942p
+  Rp1=4371.841321223
+  Cp1=4.538141294918p
+  Lp1=1.983532843425u
+  Rp2=4371.841321223
+  Cp2=4.538141294918p
+  Lp2=1.983532843425u
+  RDC1=1.60000002942979E-02
+  RDC2=1.60000002942979E-02
+  K=0.967543859162966
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874003_3.3u  1  2  3  4  PARAMS:
+  Cww=18.867p
+  Rp1=5182.94430527
+  Cp1=5.459005654292p
+  Lp1=2.658542862975u
+  Rp2=5182.94430527
+  Cp2=5.459005654292p
+  Lp2=2.658542862975u
+  RDC1=0.017750000115484
+  RDC2=0.017750000115484
+  K=0.977743431537725
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874004_4.7u  1  2  3  4  PARAMS:
+  Cww=20.012p
+  Rp1=7252.217154838
+  Cp1=4.787769338256p
+  Lp1=3.577820387445u
+  Rp2=7252.217154838
+  Cp2=4.787769338256p
+  Lp2=3.577820387445u
+  RDC1=2.14999997988343E-02
+  RDC2=2.14999997988343E-02
+  K=0.971647687479421
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874006_6.8u  1  2  3  4  PARAMS:
+  Cww=25.762p
+  Rp1=10116.401455619
+  Cp1=6.030296345694p
+  Lp1=5.819272506529u
+  Rp2=10116.401455619
+  Cp2=6.030296345694p
+  Lp2=5.819272506529u
+  RDC1=2.85000000149012E-02
+  RDC2=2.85000000149012E-02
+  K=0.967054814110566
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874101_100u  1  2  3  4  PARAMS:
+  Cww=116.482p
+  Rp1=72707.1601373
+  Cp1=8.140489777278p
+  Lp1=83.29460529805u
+  Rp2=72707.1601373
+  Cp2=8.140489777278p
+  Lp2=83.29460529805u
+  RDC1=0.261249996721745
+  RDC2=0.261249996721745
+  K=0.989836155124135
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874220_22u  1  2  3  4  PARAMS:
+  Cww=51.575p
+  Rp1=32689.83553238
+  Cp1=6.433632078578p
+  Lp1=18.75592922927u
+  Rp2=32689.83553238
+  Cp2=6.433632078578p
+  Lp2=18.75592922927u
+  RDC1=6.82500004768372E-02
+  RDC2=6.82500004768372E-02
+  K=0.983396296444086
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874470_47u  1  2  3  4  PARAMS:
+  Cww=30.316p
+  Rp1=48834.09303325
+  Cp1=6.610644800184p
+  Lp1=38.79437797437u
+  Rp2=48834.09303325
+  Cp2=6.610644800184p
+  Lp2=38.79437797437u
+  RDC1=0.127999998629093
+  RDC2=0.127999998629093
+  K=0.941562519798931
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744874100_10u  1  2  3  4  PARAMS:
+  Cww=41p
+  Rp1=15519
+  Cp1=5.485p
+  Lp1=9.558u
+  Rp2=16936
+  Cp2=5.318p
+  Lp2=10.25u
+  RDC1=0.034
+  RDC2=0.034
+  K=0.973447481891037
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1260_744871100_10u  1  2  3  4  PARAMS:
+  Cww=21p
+  Rp1=12758
+  Cp1=12.392p
+  Lp1=10.378u
+  Rp2=11256
+  Cp2=13.412p
+  Lp2=9.589u
+  RDC1=0.034
+  RDC2=0.034
+  K=0.967625960792702
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_7448700015_1.5u  1  2  3  4  PARAMS:
+  Cww=7.693p
+  Rp1=3222.084477671
+  Cp1=4.951310638861p
+  Lp1=1.27122123005u
+  Rp2=3222.084477671
+  Cp2=4.951310638861p
+  Lp2=1.27122123005u
+  RDC1=0.014750000089407
+  RDC2=0.014750000089407
+  K=0.959440559585571
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870003_3.3u  1  2  3  4  PARAMS:
+  Cww=10.87p
+  Rp1=5382.339685984
+  Cp1=7.844809681588p
+  Lp1=2.80417209167u
+  Rp2=5382.339685984
+  Cp2=7.844809681588p
+  Lp2=2.80417209167u
+  RDC1=1.89999993890524E-02
+  RDC2=1.89999993890524E-02
+  K=0.949579831963951
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870004_4.7u  1  2  3  4  PARAMS:
+  Cww=15.09p
+  Rp1=7101.347013185
+  Cp1=10.877274927613p
+  Lp1=3.612400361744u
+  Rp2=7101.347013185
+  Cp2=10.877274927613p
+  Lp2=3.612400361744u
+  RDC1=1.99999995529652E-02
+  RDC2=1.99999995529652E-02
+  K=0.961492176542446
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870006_6.8u  1  2  3  4  PARAMS:
+  Cww=18.35p
+  Rp1=10061.52839868
+  Cp1=14.121788277862p
+  Lp1=5.692951549774u
+  Rp2=10061.52839868
+  Cp2=14.121788277862p
+  Lp2=5.692951549774u
+  RDC1=2.57500004954636E-02
+  RDC2=2.57500004954636E-02
+  K=0.978478093287351
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870100_10u  1  2  3  4  PARAMS:
+  Cww=16.31p
+  Rp1=16815.56073978
+  Cp1=9.528438992978p
+  Lp1=9.326342545728u
+  Rp2=16815.56073978
+  Cp2=9.528438992978p
+  Lp2=9.326342545728u
+  RDC1=3.70000004768372E-02
+  RDC2=3.70000004768372E-02
+  K=0.954787233525386
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870101_100u  1  2  3  4  PARAMS:
+  Cww=26.86p
+  Rp1=40646.06015403
+  Cp1=35.65143913824p
+  Lp1=83.74741809743u
+  Rp2=40646.06015403
+  Cp2=35.65143913824p
+  Lp2=83.74741809743u
+  RDC1=0.217000000178814
+  RDC2=0.217000000178814
+  K=0.951572062174784
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870220_22u  1  2  3  4  PARAMS:
+  Cww=20.65p
+  Rp1=20416.76173605
+  Cp1=21.54489116668p
+  Lp1=19.66833504973u
+  Rp2=20416.76173605
+  Cp2=21.54489116668p
+  Lp2=19.66833504973u
+  RDC1=6.10000006854534E-02
+  RDC2=6.10000006854534E-02
+  K=0.959947183989084
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870221_220u  1  2  3  4  PARAMS:
+  Cww=35.47p
+  Rp1=44970.70312592
+  Cp1=48.05567458023p
+  Lp1=184.7367536363u
+  Rp2=44970.70312592
+  Cp2=48.05567458023p
+  Lp2=184.7367536363u
+  RDC1=0.452000007033348
+  RDC2=0.452000007033348
+  K=0.961599538237512
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870470_47u  1  2  3  4  PARAMS:
+  Cww=24.37p
+  Rp1=32122.07459394
+  Cp1=35.11039719801p
+  Lp1=37.88594480847u
+  Rp2=32122.07459394
+  Cp2=35.11039719801p
+  Lp2=37.88594480847u
+  RDC1=0.105750001966953
+  RDC2=0.105750001966953
+  K=0.960083064394537
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870471_470u  1  2  3  4  PARAMS:
+  Cww=39.74p
+  Rp1=58843.19082114
+  Cp1=50.91881570195p
+  Lp1=411.8554999624u
+  Rp2=58843.19082114
+  Cp2=50.91881570195p
+  Lp2=411.8554999624u
+  RDC1=0.979749977588654
+  RDC2=0.979749977588654
+  K=0.956139379483666
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870680_68u  1  2  3  4  PARAMS:
+  Cww=23.24p
+  Rp1=45061.65124881
+  Cp1=32.45509896857p
+  Lp1=57.73600099531u
+  Rp2=45061.65124881
+  Cp2=32.45509896857p
+  Lp2=57.73600099531u
+  RDC1=0.154500000178814
+  RDC2=0.154500000178814
+  K=0.940892640994621
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873001_1.5u  1  2  3  4  PARAMS:
+  Cww=11.968p
+  Rp1=3179.980596959
+  Cp1=3.69693462104p
+  Lp1=1.326037918037u
+  Rp2=3179.980596959
+  Cp2=3.69693462104p
+  Lp2=1.326037918037u
+  RDC1=1.25000001862645E-02
+  RDC2=1.25000001862645E-02
+  K=0.973492379672641
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873002_2.4u  1  2  3  4  PARAMS:
+  Cww=19.521p
+  Rp1=4235.211415115
+  Cp1=4.625030347934p
+  Lp1=1.918664789395u
+  Rp2=4235.211415115
+  Cp2=4.625030347934p
+  Lp2=1.918664789395u
+  RDC1=1.82499997317791E-02
+  RDC2=1.82499997317791E-02
+  K=0.970918155773269
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873003_3.3u  1  2  3  4  PARAMS:
+  Cww=13.548p
+  Rp1=5723.951563496
+  Cp1=5.152783352594p
+  Lp1=2.896370793236u
+  Rp2=5723.951563496
+  Cp2=5.152783352594p
+  Lp2=2.896370793236u
+  RDC1=1.70000004582107E-02
+  RDC2=1.70000004582107E-02
+  K=0.947466007467791
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873004_4.7u  1  2  3  4  PARAMS:
+  Cww=21.102p
+  Rp1=8435.054138396
+  Cp1=6.778913148162p
+  Lp1=4.571914179852u
+  Rp2=8435.054138396
+  Cp2=6.778913148162p
+  Lp2=4.571914179852u
+  RDC1=2.24999999627471E-02
+  RDC2=2.24999999627471E-02
+  K=0.949351193582894
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873100_10u  1  2  3  4  PARAMS:
+  Cww=41.216p
+  Rp1=12583.82463009
+  Cp1=10.016172539864p
+  Lp1=8.513877592868u
+  Rp2=12583.82463009
+  Cp2=10.016172539864p
+  Lp2=8.513877592868u
+  RDC1=3.54999992996454E-02
+  RDC2=3.54999992996454E-02
+  K=0.961139368819532
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873101_100u  1  2  3  4  PARAMS:
+  Cww=110.259p
+  Rp1=72334.68788369
+  Cp1=14.09239864408p
+  Lp1=82.7768210747u
+  Rp2=72334.68788369
+  Cp2=14.09239864408p
+  Lp2=82.7768210747u
+  RDC1=0.232749998569489
+  RDC2=0.232749998569489
+  K=0.98291435820526
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873150_15u  1  2  3  4  PARAMS:
+  Cww=44.002p
+  Rp1=18573.85180638
+  Cp1=10.657424319299p
+  Lp1=13.43905101848u
+  Rp2=18573.85180638
+  Cp2=10.657424319299p
+  Lp2=13.43905101848u
+  RDC1=4.42500002682209E-02
+  RDC2=4.42500002682209E-02
+  K=0.971622221204837
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873330_33u  1  2  3  4  PARAMS:
+  Cww=96.042p
+  Rp1=33295.18594266
+  Cp1=13.158260549498p
+  Lp1=29.765153975u
+  Rp2=33295.18594266
+  Cp2=13.158260549498p
+  Lp2=29.765153975u
+  RDC1=9.27499998360872E-02
+  RDC2=9.27499998360872E-02
+  K=0.991448267910977
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873470_47u  1  2  3  4  PARAMS:
+  Cww=85.902p
+  Rp1=34850.99124481
+  Cp1=12.284197732004p
+  Lp1=39.30147682288u
+  Rp2=34850.99124481
+  Cp2=12.284197732004p
+  Lp2=39.30147682288u
+  RDC1=0.105999998748302
+  RDC2=0.105999998748302
+  K=0.98720524709673
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873680_68u  1  2  3  4  PARAMS:
+  Cww=78.195p
+  Rp1=76318.8455852
+  Cp1=12.28415302188p
+  Lp1=55.18804013847u
+  Rp2=76318.8455852
+  Cp2=12.28415302188p
+  Lp2=55.18804013847u
+  RDC1=0.163499999791384
+  RDC2=0.163499999791384
+  K=0.970331864576172
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873220_22u  1  2  3  4  PARAMS:
+  Cww=138p
+  Rp1=24911
+  Cp1=9.898p
+  Lp1=19.19u
+  Rp2=25329
+  Cp2=9.434p
+  Lp2=20.139u
+  RDC1=0.051
+  RDC2=0.051
+  K=0.995215828579181
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744873221_220u  1  2  3  4  PARAMS:
+  Cww=392p
+  Rp1=76072
+  Cp1=15.289p
+  Lp1=206.26u
+  Rp2=90387
+  Cp2=14.959p
+  Lp2=210.806u
+  RDC1=0.507
+  RDC2=0.507
+  K=0.998526186664399
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870002_2.4u  1  2  3  4  PARAMS:
+  Cww=15p
+  Rp1=5225
+  Cp1=3.005p
+  Lp1=2.385u
+  Rp2=5155
+  Cp2=3.319p
+  Lp2=2.334u
+  RDC1=0.013
+  RDC2=0.013
+  K=0.921502396451939
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1280_744870151_150u  1  2  3  4  PARAMS:
+  Cww=57p
+  Rp1=44226
+  Cp1=33.023p
+  Lp1=141.066u
+  Rp2=43658
+  Cp2=34.456p
+  Lp2=135.201u
+  RDC1=0.255
+  RDC2=0.255
+  K=0.97802522121535
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878001_1.3u  1  2  3  4  PARAMS:
+  Cww=4.1875p
+  Rp1=3052.234844177
+  Cp1=4.69655033783p
+  Lp1=1.135025179597u
+  Rp2=3052.234844177
+  Cp2=4.69655033783p
+  Lp2=1.135025179597u
+  RDC1=2.67499997280538E-02
+  RDC2=2.67499997280538E-02
+  K=0.960317459801232
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878002_2.4u  1  2  3  4  PARAMS:
+  Cww=4.9625p
+  Rp1=5302.644154298
+  Cp1=4.396748958066p
+  Lp1=2.14408628271u
+  Rp2=5302.644154298
+  Cp2=4.396748958066p
+  Lp2=2.14408628271u
+  RDC1=4.05000001192093E-02
+  RDC2=4.05000001192093E-02
+  K=0.941544882014607
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878003_3.3u  1  2  3  4  PARAMS:
+  Cww=4.13p
+  Rp1=6277.400426277
+  Cp1=4.327343439359p
+  Lp1=2.829370009363u
+  Rp2=6277.400426277
+  Cp2=4.327343439359p
+  Lp2=2.829370009363u
+  RDC1=4.55000000074506E-02
+  RDC2=4.55000000074506E-02
+  K=0.94551281906777
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878004_4.7u  1  2  3  4  PARAMS:
+  Cww=4.92p
+  Rp1=8272.09663569
+  Cp1=5.400933342016p
+  Lp1=3.923743823943u
+  Rp2=8272.09663569
+  Cp2=5.400933342016p
+  Lp2=3.923743823943u
+  RDC1=6.32500005885959E-02
+  RDC2=6.32500005885959E-02
+  K=0.908994710922295
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878005_5.6u  1  2  3  4  PARAMS:
+  Cww=4.53p
+  Rp1=9428.694075054
+  Cp1=6.074558702798p
+  Lp1=5.336219581368u
+  Rp2=9428.694075054
+  Cp2=6.074558702798p
+  Lp2=5.336219581368u
+  RDC1=8.37500002235174E-02
+  RDC2=8.37500002235174E-02
+  K=0.919672132166314
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878006_6.8u  1  2  3  4  PARAMS:
+  Cww=4.95p
+  Rp1=11220.88323414
+  Cp1=6.088135735101p
+  Lp1=6.117137346139u
+  Rp2=11220.88323414
+  Cp2=6.088135735101p
+  Lp2=6.117137346139u
+  RDC1=8.95000025629997E-02
+  RDC2=8.95000025629997E-02
+  K=0.921795797899602
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878008_8.2u  1  2  3  4  PARAMS:
+  Cww=5.305p
+  Rp1=11772.616750928
+  Cp1=6.316033400206p
+  Lp1=6.925907479861u
+  Rp2=11772.616750928
+  Cp2=6.316033400206p
+  Lp2=6.925907479861u
+  RDC1=0.103250002488494
+  RDC2=0.103250002488494
+  K=0.915596330074557
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878100_10u  1  2  3  4  PARAMS:
+  Cww=5.35p
+  Rp1=14085.14549534
+  Cp1=5.803172523208p
+  Lp1=8.442790496906u
+  Rp2=14085.14549534
+  Cp2=5.803172523208p
+  Lp2=8.442790496906u
+  RDC1=0.127750001847744
+  RDC2=0.127750001847744
+  K=0.922675024972665
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878101_100u  1  2  3  4  PARAMS:
+  Cww=9.41p
+  Rp1=63426.1945521
+  Cp1=10.419700222087p
+  Lp1=87.02321671935u
+  Rp2=63426.1945521
+  Cp2=10.419700222087p
+  Lp2=87.02321671935u
+  RDC1=1.16899999976158
+  RDC2=1.16899999976158
+  K=0.938248462535577
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878220_22u  1  2  3  4  PARAMS:
+  Cww=6.51p
+  Rp1=23974.33598126
+  Cp1=7.743012783924p
+  Lp1=18.67164732777u
+  Rp2=23974.33598126
+  Cp2=7.743012783924p
+  Lp2=18.67164732777u
+  RDC1=0.244000002741814
+  RDC2=0.244000002741814
+  K=0.918906395956803
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7332_744878470_47u  1  2  3  4  PARAMS:
+  Cww=9.525p
+  Rp1=39039.49084463
+  Cp1=9.373403111728p
+  Lp1=43.44145091395u
+  Rp2=39039.49084463
+  Cp2=9.373403111728p
+  Lp2=43.44145091395u
+  RDC1=0.569999992847443
+  RDC2=0.569999992847443
+  K=0.944001678058741
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877001_1.8u  1  2  3  4  PARAMS:
+  Cww=4.94p
+  Rp1=3735.482360635
+  Cp1=4.157668652089p
+  Lp1=1.483081091204u
+  Rp2=3735.482360635
+  Cp2=4.157668652089p
+  Lp2=1.483081091204u
+  RDC1=0.02625000057742
+  RDC2=0.02625000057742
+  K=0.968553458367985
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877002_2.4u  1  2  3  4  PARAMS:
+  Cww=6.35p
+  Rp1=4399.661140784
+  Cp1=5.306931952009p
+  Lp1=2.031508130452u
+  Rp2=4399.661140784
+  Cp2=5.306931952009p
+  Lp2=2.031508130452u
+  RDC1=3.05000012740493E-02
+  RDC2=3.05000012740493E-02
+  K=0.912499999006589
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877003_3.3u  1  2  3  4  PARAMS:
+  Cww=7.75p
+  Rp1=6729.932531648
+  Cp1=6.276574117184p
+  Lp1=3.24681399793u
+  Rp2=6729.932531648
+  Cp2=6.276574117184p
+  Lp2=3.24681399793u
+  RDC1=4.17499989271164E-02
+  RDC2=4.17499989271164E-02
+  K=0.955801103257612
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877004_4.7u  1  2  3  4  PARAMS:
+  Cww=6.75p
+  Rp1=7330.545982911
+  Cp1=6.625178973507p
+  Lp1=3.800255270261u
+  Rp2=7330.545982911
+  Cp2=6.625178973507p
+  Lp2=3.800255270261u
+  RDC1=4.62500005960464E-02
+  RDC2=4.62500005960464E-02
+  K=0.935267854600727
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877005_5.6u  1  2  3  4  PARAMS:
+  Cww=6.645p
+  Rp1=9678.501698923
+  Cp1=5.246342504626p
+  Lp1=4.815919780821u
+  Rp2=9678.501698923
+  Cp2=5.246342504626p
+  Lp2=4.815919780821u
+  RDC1=6.64999997243285E-02
+  RDC2=6.64999997243285E-02
+  K=0.938125567833223
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877006_6.8u  1  2  3  4  PARAMS:
+  Cww=7.1625p
+  Rp1=11623.77221658
+  Cp1=7.115754050699p
+  Lp1=6.536803658278u
+  Rp2=11623.77221658
+  Cp2=7.115754050699p
+  Lp2=6.536803658278u
+  RDC1=7.87499994039536E-02
+  RDC2=7.87499994039536E-02
+  K=0.946575341975852
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877008_8.2u  1  2  3  4  PARAMS:
+  Cww=8.2p
+  Rp1=12142.64744534
+  Cp1=7.866482393082p
+  Lp1=7.874363281789u
+  Rp2=12142.64744534
+  Cp2=7.866482393082p
+  Lp2=7.874363281789u
+  RDC1=8.32500010728836E-02
+  RDC2=8.32500010728836E-02
+  K=0.960045662954863
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877100_10u  1  2  3  4  PARAMS:
+  Cww=8.415p
+  Rp1=11554.12199734
+  Cp1=10.971494144547p
+  Lp1=8.504394301672u
+  Rp2=11554.12199734
+  Cp2=10.971494144547p
+  Lp2=8.504394301672u
+  RDC1=8.99999998509884E-02
+  RDC2=8.99999998509884E-02
+  K=0.947530863334485
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877101_100u  1  2  3  4  PARAMS:
+  Cww=13.17p
+  Rp1=60156.7589142
+  Cp1=16.66620330062p
+  Lp1=89.00392736262u
+  Rp2=60156.7589142
+  Cp2=16.66620330062p
+  Lp2=89.00392736262u
+  RDC1=0.901500016450881
+  RDC2=0.901500016450881
+  K=0.957361554101469
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877220_22u  1  2  3  4  PARAMS:
+  Cww=10.37p
+  Rp1=20724.9180642
+  Cp1=12.8132294158889p
+  Lp1=19.3530956566778u
+  Rp2=20724.9180642
+  Cp2=12.8132294158889p
+  Lp2=19.3530956566778u
+  RDC1=0.190500002354383
+  RDC2=0.190500002354383
+  K=0.956810631447276
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 7345_744877330_33u  1  2  3  4  PARAMS:
+  Cww=9.715p
+  Rp1=30858.1675609
+  Cp1=11.079332484208p
+  Lp1=30.58837073111u
+  Rp2=30858.1675609
+  Cp2=11.079332484208p
+  Lp2=30.58837073111u
+  RDC1=0.338250003755093
+  RDC2=0.338250003755093
+  K=0.934893489056838
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
