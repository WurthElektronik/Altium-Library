**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Film Capacitor
* Matchcode:             WCAP-FTDB
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         7/11/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 890484427001CS_35uF 1 2
Rser 1 3 0.0058
Lser 2 4 0.0000000158
C1 3 4 0.000035
Rpar 3 4 2000000000
.ends 890484427001CS_35uF
*******
.subckt 890484428002CS_1uF 1 2
Rser 1 3 0.0495
Lser 2 4 0.0000000135
C1 3 4 0.000001
Rpar 3 4 285714286
.ends 890484428002CS_1uF
*******
.subckt 890484429001CS_50uF 1 2
Rser 1 3 0.00655
Lser 2 4 0.0000000479
C1 3 4 0.00005
Rpar 3 4 133333333
.ends 890484429001CS_50uF
*******
.subckt 890494427003CS_3uF 1 2
Rser 1 3 0.021
Lser 2 4 0.0000000173
C1 3 4 0.000003
Rpar 3 4 3333333333
.ends 890494427003CS_3uF
*******
.subckt 890494428004CS_3uF 1 2
Rser 1 3 0.02
Lser 2 4 0.0000000153
C1 3 4 0.000003
Rpar 3 4 400000000
.ends 890494428004CS_3uF
*******
.subckt 890494429003CS_25uF 1 2
Rser 1 3 0.00725
Lser 2 4 0.0000000325
C1 3 4 0.000025
Rpar 3 4 250000000
.ends 890494429003CS_25uF
*******
.subckt 890494429005CS_10uF 1 2
Rser 1 3 0.013
Lser 2 4 0.0000000133
C1 3 4 0.00001
Rpar 3 4 200000000
.ends 890494429005CS_10uF
*******
.subckt 890714429003CS_10uF 1 2
Rser 1 3 0.014
Lser 2 4 0.00000003
C1 3 4 0.00001
Rpar 3 4 200000000
.ends 890714429003CS_10uF
*******
.subckt 890724427001CS_5uF 1 2
Rser 1 3 0.017
Lser 2 4 0.0000000122
C1 3 4 0.000005
Rpar 3 4 10000000000
.ends 890724427001CS_5uF
*******
.subckt 890724427010CS_10uF 1 2
Rser 1 3 0.0115
Lser 2 4 0.0000000134
C1 3 4 0.00001
Rpar 3 4 1000000000
.ends 890724427010CS_10uF
*******
.subckt 890724429005CS_25uF 1 2
Rser 1 3 0.0075
Lser 2 4 0.0000000349
C1 3 4 0.000025
Rpar 3 4 200000000
.ends 890724429005CS_25uF
*******
.subckt 890724429010CS_1uF 1 2
Rser 1 3 0.05
Lser 2 4 0.0000000114
C1 3 4 0.000001
Rpar 3 4 133333333
.ends 890724429010CS_1uF
*******
.subckt 890734427005CS_25uF 1 2
Rser 1 3 0.007
Lser 2 4 0.0000000287
C1 3 4 0.000025
Rpar 3 4 3333333333
.ends 890734427005CS_25uF
*******
.subckt 890734428004CS_50uF 1 2
Rser 1 3 0.006
Lser 2 4 0.0000000284
C1 3 4 0.00005
Rpar 3 4 666666667
.ends 890734428004CS_50uF
*******
.subckt 890734428008CS_15uF 1 2
Rser 1 3 0.0105
Lser 2 4 0.0000000321
C1 3 4 0.000015
Rpar 3 4 333333333
.ends 890734428008CS_15uF
*******
.subckt 890734429007CS_40uF 1 2
Rser 1 3 0.0047
Lser 2 4 0.0000000228
C1 3 4 0.00004
Rpar 3 4 200000000
.ends 890734429007CS_40uF
*******
.subckt 890744427001CS_75uF 1 2
Rser 1 3 0.00614
Lser 2 4 0.0000000263
C1 3 4 0.000075
Rpar 3 4 10000000000
.ends 890744427001CS_75uF
*******
.subckt 890744427005CS_50uF 1 2
Rser 1 3 0.006
Lser 2 4 0.0000000272
C1 3 4 0.00005
Rpar 3 4 2000000000
.ends 890744427005CS_50uF
*******
.subckt 890744428006CS_30uF 1 2
Rser 1 3 0.00605
Lser 2 4 0.0000000369
C1 3 4 0.00003
Rpar 3 4 400000000
.ends 890744428006CS_30uF
*******
.subckt 890744429002CS_40uF 1 2
Rser 1 3 0.00572
Lser 2 4 0.0000000443
C1 3 4 0.00004
Rpar 3 4 400000000
.ends 890744429002CS_40uF
*******
.subckt 890744429005CS_60uF 1 2
Rser 1 3 0.00585
Lser 2 4 0.0000000252
C1 3 4 0.00006
Rpar 3 4 250000000
.ends 890744429005CS_60uF
*******
.subckt 890764427009CS_40uF 1 2
Rser 1 3 0.00824
Lser 2 4 0.0000000294
C1 3 4 0.00004
Rpar 3 4 1000000000
.ends 890764427009CS_40uF
*******
.subckt 890764428004CS_75uF 1 2
Rser 1 3 0.004
Lser 2 4 0.000000032
C1 3 4 0.000075
Rpar 3 4 250000000
.ends 890764428004CS_75uF
*******
.subckt 890764429002CS_5uF 1 2
Rser 1 3 0.016
Lser 2 4 0.0000000155
C1 3 4 0.000005
Rpar 3 4 166666667
.ends 890764429002CS_5uF
*******
