**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT High Current Inductor
* Matchcode:              WE-HCF 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-09
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 2013_7443630070_0.7u 1 2
Rp 1 2 280.93
Cp 1 2 5.973p
Rs 1 N3 0.000829
L1 N3 2 0.667811u
.ends 2013_7443630070_0.7u
*******
.subckt 2013_7443630140_1.4u 1 2
Rp 1 2 525.687
Cp 1 2 5.479p
Rs 1 N3 0.001083
L1 N3 2 1.307u
.ends 2013_7443630140_1.4u
*******
.subckt 2013_7443630220_2.2u 1 2
Rp 1 2 830.152
Cp 1 2 5.727p
Rs 1 N3 0.0015
L1 N3 2 1.995u
.ends 2013_7443630220_2.2u
*******
.subckt 2013_7443630310_3.1u 1 2
Rp 1 2 1379
Cp 1 2 7.104p
Rs 1 N3 0.002085
L1 N3 2 2.887u
.ends 2013_7443630310_3.1u
*******
.subckt 2013_7443630420_4.2u 1 2
Rp 1 2 1709
Cp 1 2 5.527p
Rs 1 N3 0.003038
L1 N3 2 3.71u
.ends 2013_7443630420_4.2u
*******
.subckt 2013_7443630550_5.5u 1 2
Rp 1 2 2374
Cp 1 2 5.469p
Rs 1 N3 0.004
L1 N3 2 5.777u
.ends 2013_7443630550_5.5u
*******
.subckt 2013_7443630700_7u 1 2
Rp 1 2 3136
Cp 1 2 5.159p
Rs 1 N3 0.005608
L1 N3 2 6.346u
.ends 2013_7443630700_7u
*******
.subckt 2013_7443630860_8.6u 1 2
Rp 1 2 3955
Cp 1 2 5.388p
Rs 1 N3 0.007186
L1 N3 2 7.677u
.ends 2013_7443630860_8.6u
*******
.subckt 2013_7443631000_10u 1 2
Rp 1 2 4405
Cp 1 2 4.764p
Rs 1 N3 0.00796
L1 N3 2 8.683u
.ends 2013_7443631000_10u
*******
.subckt 2013_7443631500_15u 1 2
Rp 1 2 6395
Cp 1 2 6.255p
Rs 1 N3 0.0087
L1 N3 2 13.341u
.ends 2013_7443631500_15u
*******
.subckt 2013_7443632200_22u 1 2
Rp 1 2 8040
Cp 1 2 5.208p
Rs 1 N3 0.01065
L1 N3 2 20.243u
.ends 2013_7443632200_22u
*******
.subckt 2013_7443633300_33u 1 2
Rp 1 2 8318
Cp 1 2 6.362p
Rs 1 N3 0.0114
L1 N3 2 31.744u
.ends 2013_7443633300_33u
*******
.subckt 2013_7443634700_47u 1 2
Rp 1 2 11320
Cp 1 2 7.067p
Rs 1 N3 0.0122
L1 N3 2 42.742u
.ends 2013_7443634700_47u
*******
.subckt 2815_74436410150_1.5u 1 2
Rp 1 2 1082
Cp 1 2 9.173p
Rs 1 N3 0.00133
L1 N3 2 1.486u
.ends 2815_74436410150_1.5u
*******
.subckt 2815_74436410220_2.2u 1 2
Rp 1 2 1034
Cp 1 2 10.39p
Rs 1 N3 0.00133
L1 N3 2 2.273u
.ends 2815_74436410220_2.2u
*******
.subckt 2815_74436410330_3.3u 1 2
Rp 1 2 1179
Cp 1 2 11.15p
Rs 1 N3 0.00133
L1 N3 2 3.26u
.ends 2815_74436410330_3.3u
*******
.subckt 2815_74436410470_4.7u 1 2
Rp 1 2 1219
Cp 1 2 12.36p
Rs 1 N3 0.00133
L1 N3 2 4.45u
.ends 2815_74436410470_4.7u
*******
.subckt 2815_74436410680_6.8u 1 2
Rp 1 2 1214
Cp 1 2 13.33p
Rs 1 N3 0.00133
L1 N3 2 6.56u
.ends 2815_74436410680_6.8u
*******
.subckt 2815_74436411000_10u 1 2
Rp 1 2 1230
Cp 1 2 13.79p
Rs 1 N3 0.00133
L1 N3 2 10.02u
.ends 2815_74436411000_10u
*******
.subckt 2815_74436411500_15u 1 2
Rp 1 2 1294
Cp 1 2 14.97p
Rs 1 N3 0.00133
L1 N3 2 14.78u
.ends 2815_74436411500_15u
*******
.subckt 2815_74436412200_22u 1 2
Rp 1 2 1395
Cp 1 2 17.1p
Rs 1 N3 0.00133
L1 N3 2 22.83u
.ends 2815_74436412200_22u
*******
.subckt 2815_74436413300_33u 1 2
Rp 1 2 1543
Cp 1 2 18.36p
Rs 1 N3 0.00133
L1 N3 2 35.15u
.ends 2815_74436413300_33u
*******
.subckt 2818_7443640330_3.3u 1 2
Rp 1 2 1120
Cp 1 2 17.55p
Rs 1 N3 0.0024
L1 N3 2 3.3u
.ends 2818_7443640330_3.3u
*******
.subckt 2818_7443640470_4.7u 1 2
Rp 1 2 1190
Cp 1 2 17.91p
Rs 1 N3 0.0024
L1 N3 2 4.7u
.ends 2818_7443640470_4.7u
*******
.subckt 2818_7443640680_6.8u 1 2
Rp 1 2 1230
Cp 1 2 18.73p
Rs 1 N3 0.0024
L1 N3 2 6.8u
.ends 2818_7443640680_6.8u
*******
.subckt 2818_7443641000_10u 1 2
Rp 1 2 1310
Cp 1 2 18.05p
Rs 1 N3 0.0024
L1 N3 2 10u
.ends 2818_7443641000_10u
*******
.subckt 2818_7443641500_15u 1 2
Rp 1 2 1330
Cp 1 2 18.29p
Rs 1 N3 0.0024
L1 N3 2 15u
.ends 2818_7443641500_15u
*******
.subckt 2818_7443642200_22u 1 2
Rp 1 2 1440
Cp 1 2 19.93p
Rs 1 N3 0.0024
L1 N3 2 22u
.ends 2818_7443642200_22u
*******
.subckt 2818_7443643300_33u 1 2
Rp 1 2 1470
Cp 1 2 17.8p
Rs 1 N3 0.0024
L1 N3 2 33u
.ends 2818_7443643300_33u
*******
.subckt 2818B_7443640100B_1u 1 2
Rp 1 2 389.52
Cp 1 2 4.73958514312p
Rs 1 N3 0.00044
L1 N3 2 1.06469752848u
.ends 2818B_7443640100B_1u
*******
.subckt 2818B_7443640150B_1.5u 1 2
Rp 1 2 422.7
Cp 1 2 6.60175663697p
Rs 1 N3 0.00044
L1 N3 2 1.72246545684u
.ends 2818B_7443640150B_1.5u
*******
.subckt 2818B_7443640330B_3.3u 1 2
Rp 1 2 1113
Cp 1 2 8.386p
Rs 1 N3 0.00044
L1 N3 2 3.374u
.ends 2818B_7443640330B_3.3u
*******
.subckt 2818B_7443640470B_4.7u 1 2
Rp 1 2 1213
Cp 1 2 9.419p
Rs 1 N3 0.00044
L1 N3 2 4.856u
.ends 2818B_7443640470B_4.7u
*******
.subckt 2818B_7443640680B_6.8u 1 2
Rp 1 2 1121
Cp 1 2 11.063p
Rs 1 N3 0.00044
L1 N3 2 6.45u
.ends 2818B_7443640680B_6.8u
*******
.subckt 2818B_7443641000B_10u 1 2
Rp 1 2 1140
Cp 1 2 12.35p
Rs 1 N3 0.00044
L1 N3 2 9.034u
.ends 2818B_7443641000B_10u
*******
.subckt 2920_74437429203101_100u 1 2
Rp 1 2 18328
Cp 1 2 13.548p
Rs 1 N3 0.0359
L1 N3 2 104.807u
.ends 2920_74437429203101_100u
*******
.subckt 2920_74437429203151_150u 1 2
Rp 1 2 23820
Cp 1 2 12.272p
Rs 1 N3 0.03885
L1 N3 2 141.778u
.ends 2920_74437429203151_150u
*******
.subckt 2920_74437429203330_33u 1 2
Rp 1 2 6230
Cp 1 2 11.191p
Rs 1 N3 0.0153
L1 N3 2 32.98u
.ends 2920_74437429203330_33u
*******
.subckt 2920_74437429203470_47u 1 2
Rp 1 2 9270
Cp 1 2 8.882p
Rs 1 N3 0.0193
L1 N3 2 48.005u
.ends 2920_74437429203470_47u
*******
.subckt 2920_74437429203680_68u 1 2
Rp 1 2 10735
Cp 1 2 12.705p
Rs 1 N3 0.0222
L1 N3 2 70.591u
.ends 2920_74437429203680_68u
*******
.subckt 2920_74437529203101_100u 1 2
Rp 1 2 21321
Cp 1 2 13.609p
Rs 1 N3 0.0229
L1 N3 2 104.516u
.ends 2920_74437529203101_100u
*******
.subckt 2920_74437529203151_150u 1 2
Rp 1 2 35180
Cp 1 2 13.607p
Rs 1 N3 0.0306
L1 N3 2 176.178u
.ends 2920_74437529203151_150u
*******
.subckt 2920_74437529203220_22u 1 2
Rp 1 2 4184
Cp 1 2 12.758p
Rs 1 N3 0.0049
L1 N3 2 22.743u
.ends 2920_74437529203220_22u
*******
.subckt 2920_74437529203221_220u 1 2
Rp 1 2 35623
Cp 1 2 14.233p
Rs 1 N3 0.03645
L1 N3 2 213.326u
.ends 2920_74437529203221_220u
*******
.subckt 2920_74437529203330_33u 1 2
Rp 1 2 5743
Cp 1 2 14.457p
Rs 1 N3 0.0069
L1 N3 2 32.553u
.ends 2920_74437529203330_33u
*******
.subckt 2920_74437529203331_330u 1 2
Rp 1 2 58482
Cp 1 2 13.251p
Rs 1 N3 0.07045
L1 N3 2 347.127u
.ends 2920_74437529203331_330u
*******
.subckt 2920_74437529203470_47u 1 2
Rp 1 2 7147
Cp 1 2 11.864p
Rs 1 N3 0.0088
L1 N3 2 47.09u
.ends 2920_74437529203470_47u
*******
.subckt 2920_74437529203471_470u 1 2
Rp 1 2 78896
Cp 1 2 19.022p
Rs 1 N3 0.08345
L1 N3 2 455.031u
.ends 2920_74437529203471_470u
*******
.subckt 2920_74437529203680_68u 1 2
Rp 1 2 11503
Cp 1 2 12.335p
Rs 1 N3 0.0103
L1 N3 2 64.695u
.ends 2920_74437529203680_68u
*******
.subckt 2920_74437529203681_680u 1 2
Rp 1 2 85440
Cp 1 2 22.797p
Rs 1 N3 0.1183
L1 N3 2 867.917u
.ends 2920_74437529203681_680u
*******
.subckt 2010_7443642010100_1u 1 2
Rp 1 2 265.601
Cp 1 2 13.505p
Rs 1 N3 0.84m
L1 N3 2 927.701n
.ends 2010_7443642010100_1u
*******
.subckt 2010_7443642010120_1.2u 1 2
Rp 1 2 271.844
Cp 1 2 13.069p
Rs 1 N3 0.84m
L1 N3 2 1.079u
.ends 2010_7443642010120_1.2u
*******
.subckt 2010_7443642010200_2u 1 2
Rp 1 2 308.651
Cp 1 2 16.021p
Rs 1 N3 0.84m
L1 N3 2 1.749u
.ends 2010_7443642010200_2u
*******