**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Dual Powerchoke 
* Matchcode:              WE-DPC 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 5838_7448844010_1u  1  2  3  4  PARAMS:
+  Cww=6.2p
+  Rp1=429
+  Cp1=2.58p
+  Lp1=1.031u
+  Rp2=457
+  Cp2=2.361p
+  Lp2=1.127u
+  RDC1=0.017
+  RDC2=0.017
+  K=0.91214034007931
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844022_2.2u  1  2  3  4  PARAMS:
+  Cww=9.8p
+  Rp1=1461
+  Cp1=2.822p
+  Lp1=2.162u
+  Rp2=1446
+  Cp2=2.333p
+  Lp2=2.114u
+  RDC1=0.028
+  RDC2=0.028
+  K=0.960113629638795
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844033_3.3u  1  2  3  4  PARAMS:
+  Cww=12p
+  Rp1=2267
+  Cp1=3.321p
+  Lp1=3.307u
+  Rp2=2260
+  Cp2=3.305p
+  Lp2=3.382u
+  RDC1=0.034
+  RDC2=0.034
+  K=0.971253485622231
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844047_4.7u  1  2  3  4  PARAMS:
+  Cww=14p
+  Rp1=3591
+  Cp1=3.123p
+  Lp1=5.309u
+  Rp2=3588
+  Cp2=3.114p
+  Lp2=5.324u
+  RDC1=0.047
+  RDC2=0.047
+  K=0.979035565389671
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844068_6.8u  1  2  3  4  PARAMS:
+  Cww=16p
+  Rp1=5036
+  Cp1=3.513p
+  Lp1=7.215u
+  Rp2=4915
+  Cp2=3.412p
+  Lp2=7.301u
+  RDC1=0.058
+  RDC2=0.058
+  K=0.982942760585903
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844100_10u  1  2  3  4  PARAMS:
+  Cww=18p
+  Rp1=6481
+  Cp1=3.658p
+  Lp1=10.064u
+  Rp2=6790
+  Cp2=3.637p
+  Lp2=10.122u
+  RDC1=0.08
+  RDC2=0.08
+  K=0.987319603775799
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844150_15u  1  2  3  4  PARAMS:
+  Cww=26p
+  Rp1=9883
+  Cp1=3.112p
+  Lp1=15.297u
+  Rp2=9817
+  Cp2=3.1p
+  Lp2=15.487u
+  RDC1=0.13
+  RDC2=0.13
+  K=0.990689995239008
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844220_22u  1  2  3  4  PARAMS:
+  Cww=37p
+  Rp1=13155
+  Cp1=3.458p
+  Lp1=19.733u
+  Rp2=13014
+  Cp2=3.444p
+  Lp2=19.816u
+  RDC1=0.169
+  RDC2=0.169
+  K=0.992013562957135
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844330_33u  1  2  3  4  PARAMS:
+  Cww=40p
+  Rp1=20313
+  Cp1=3.751p
+  Lp1=33.361u
+  Rp2=21415
+  Cp2=3.704p
+  Lp2=33.15u
+  RDC1=0.22
+  RDC2=0.22
+  K=0.992883770548286
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 5838_7448844470_47u  1  2  3  4  PARAMS:
+  Cww=47p
+  Rp1=27605
+  Cp1=3.898p
+  Lp1=43.106u
+  Rp2=26311
+  Cp2=3.843p
+  Lp2=44.746u
+  RDC1=0.24
+  RDC2=0.24
+  K=0.993596518992086
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
