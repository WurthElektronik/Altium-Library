**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT High Current Flat Wire Inductor 
* Matchcode:              WE-HCM 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-09
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1050_744303012_0.12u  1 2
Rp 1 2 71.54
Cp 1 2 11p
Rs 1 N3 0.000325
L1 N3 2 0.12144u
.ends 1050_744303012_0.12u 
*******
.subckt 1050_744303015_0.155u  1 2
Rp 1 2 69.77
Cp 1 2 20.21p
Rs 1 N3 0.000325
L1 N3 2 0.1706u
.ends 1050_744303015_0.155u 
*******
.subckt 1050_744303022_0.22u  1 2
Rp 1 2 84.88
Cp 1 2 18.52p
Rs 1 N3 0.000325
L1 N3 2 0.26084u
.ends 1050_744303022_0.22u 
*******
.subckt 1052_744306020_0.2u  1 2
Rp 1 2 53.9
Cp 1 2 0.927p
Rs 1 N3 0.0003
L1 N3 2 0.22133u
.ends 1052_744306020_0.2u 
*******
.subckt 1052_744306025_0.25u  1 2
Rp 1 2 55.47
Cp 1 2 0.526p
Rs 1 N3 0.0003
L1 N3 2 0.32579u
.ends 1052_744306025_0.25u 
*******
.subckt 1052_744306030_0.3u  1 2
Rp 1 2 53.22
Cp 1 2 29.61p
Rs 1 N3 0.0003
L1 N3 2 0.36692u
.ends 1052_744306030_0.3u 
*******
.subckt 1070_744308015_0.15u  1 2
Rp 1 2 57.41
Cp 1 2 1.9p
Rs 1 N3 0.00037
L1 N3 2 0.19782u
.ends 1070_744308015_0.15u 
*******
.subckt 1070_744308020_0.2u  1 2
Rp 1 2 61.66
Cp 1 2 1.327p
Rs 1 N3 0.00037
L1 N3 2 0.21483u
.ends 1070_744308020_0.2u 
*******
.subckt 1070_744308025_0.25u  1 2
Rp 1 2 64.55
Cp 1 2 1.694p
Rs 1 N3 0.00037
L1 N3 2 0.29257u
.ends 1070_744308025_0.25u 
*******
.subckt 1070_744308033_0.33u  1 2
Rp 1 2 69.73
Cp 1 2 0.991p
Rs 1 N3 0.00037
L1 N3 2 0.38974u
.ends 1070_744308033_0.33u 
*******
.subckt 1070_744308040_0.4u  1 2
Rp 1 2 50.667
Cp 1 2 21.667p
Rs 1 N3 0.00037
L1 N3 2 0.501667u
.ends 1070_744308040_0.4u 
*******
.subckt 1190_744301025_0.25u  1 2
Rp 1 2 45.7
Cp 1 2 1.13p
Rs 1 N3 0.00032
L1 N3 2 0.281u
.ends 1190_744301025_0.25u 
*******
.subckt 1190_744301033_0.33u  1 2
Rp 1 2 34.58
Cp 1 2 7.25p
Rs 1 N3 0.00032
L1 N3 2 0.284u
.ends 1190_744301033_0.33u 
*******
.subckt 1190_744301047_0.47u  1 2
Rp 1 2 47.76
Cp 1 2 0.1283p
Rs 1 N3 0.00032
L1 N3 2 0.486u
.ends 1190_744301047_0.47u 
*******
.subckt 1240_744304010_0.1u  1 2
Rp 1 2 41.01
Cp 1 2 9.08p
Rs 1 N3 0.00017
L1 N3 2 0.1065u
.ends 1240_744304010_0.1u 
*******
.subckt 1240_744304016_0.16u  1 2
Rp 1 2 59.08
Cp 1 2 17.7p
Rs 1 N3 0.00017
L1 N3 2 0.1722u
.ends 1240_744304016_0.16u 
*******
.subckt 1240_744304022_0.22u  1 2
Rp 1 2 51.23
Cp 1 2 22.68p
Rs 1 N3 0.00017
L1 N3 2 0.223u
.ends 1240_744304022_0.22u 
*******
.subckt 1350_744305022_0.22u  1 2
Rp 1 2 55.28
Cp 1 2 0.247p
Rs 1 N3 0.000155
L1 N3 2 0.29797u
.ends 1350_744305022_0.22u 
*******
.subckt 1350_744305033_0.33u  1 2
Rp 1 2 58.24
Cp 1 2 40.74p
Rs 1 N3 0.000155
L1 N3 2 0.36362u
.ends 1350_744305033_0.33u 
*******
.subckt 1350_744305040_0.4u  1 2
Rp 1 2 62.85
Cp 1 2 22.58p
Rs 1 N3 0.000155
L1 N3 2 0.48324u
.ends 1350_744305040_0.4u 
*******
.subckt 1390_744309012_0.12u  1 2
Rp 1 2 41
Cp 1 2 26p
Rs 1 N3 0.000165
L1 N3 2 0.12u
.ends 1390_744309012_0.12u 
*******
.subckt 1390_744309025_0.25u  1 2
Rp 1 2 41.08
Cp 1 2 0.994p
Rs 1 N3 0.000165
L1 N3 2 0.283u
.ends 1390_744309025_0.25u 
*******
.subckt 1390_744309033_0.33u  1 2
Rp 1 2 41.5
Cp 1 2 2.38p
Rs 1 N3 0.000165
L1 N3 2 0.392u
.ends 1390_744309033_0.33u 
*******
.subckt 1390_744309047_0.47u  1 2
Rp 1 2 39.42
Cp 1 2 4.62p
Rs 1 N3 0.000165
L1 N3 2 0.599u
.ends 1390_744309047_0.47u 
*******
.subckt 7050_744302007_0.072u  1 2
Rp 1 2 42.42
Cp 1 2 18.39p
Rs 1 N3 0.000235
L1 N3 2 0.077366u
.ends 7050_744302007_0.072u 
*******
.subckt 7050_744302010_0.105u  1 2
Rp 1 2 35.46
Cp 1 2 50.45p
Rs 1 N3 0.000235
L1 N3 2 0.1178u
.ends 7050_744302010_0.105u 
*******
.subckt 7050_744302015_0.15u  1 2
Rp 1 2 51.16
Cp 1 2 46.07p
Rs 1 N3 0.000235
L1 N3 2 0.16722u
.ends 7050_744302015_0.15u 
*******
.subckt 7070_744307012_0.12u  1 2
Rp 1 2 41.79
Cp 1 2 0.694p
Rs 1 N3 0.00033
L1 N3 2 0.16394u
.ends 7070_744307012_0.12u 
*******
.subckt 7070_744307016_0.16u  1 2
Rp 1 2 42.31
Cp 1 2 0.4289p
Rs 1 N3 0.00033
L1 N3 2 0.18954u
.ends 7070_744307016_0.16u 
*******
.subckt 7070_744307022_0.22u  1 2
Rp 1 2 47.3
Cp 1 2 0.664p
Rs 1 N3 0.00033
L1 N3 2 0.2489u
.ends 7070_744307022_0.22u 
*******
.subckt 1078_7443081010_0.1u  1 2
Rp 1 2 36.968
Cp 1 2 300.126p
Rs 1 N3 0.00029
L1 N3 2 0.1u
.ends 1078_7443081010_0.1u 
*******
.subckt 1078_7443081012_0.12u  1 2
Rp 1 2 36.968
Cp 1 2 353.854p
Rs 1 N3 0.00029
L1 N3 2 0.12u
.ends 1078_7443081012_0.12u 
*******
.subckt 1078_7443081015_0.15u  1 2
Rp 1 2 37.033
Cp 1 2 31.354p
Rs 1 N3 0.00029
L1 N3 2 0.15u
.ends 1078_7443081015_0.15u 
*******
.subckt 1078_7443081018_0.18u  1 2
Rp 1 2 38.971
Cp 1 2 690.847p
Rs 1 N3 0.00029
L1 N3 2 0.18u
.ends 1078_7443081018_0.18u 
*******
.subckt 1078_7443081022_0.22u  1 2
Rp 1 2 42.567
Cp 1 2 1.075p
Rs 1 N3 0.00029
L1 N3 2 0.22u
.ends 1078_7443081022_0.22u 
*******
.subckt 1078_7443081030_0.3u  1 2
Rp 1 2 43.708
Cp 1 2 1.692p
Rs 1 N3 0.00029
L1 N3 2 0.3u
.ends 1078_7443081030_0.3u 
*******
.subckt 1078_7443081040_0.4u  1 2
Rp 1 2 48.258
Cp 1 2 2.687p
Rs 1 N3 0.00029
L1 N3 2 0.4u
.ends 1078_7443081040_0.4u 
*******
.subckt 1088_7443082010_0.1u  1 2
Rp 1 2 30.8
Cp 1 2 30.47p
Rs 1 N3 0.00018
L1 N3 2 0.1002u
.ends 1088_7443082010_0.1u 
*******
.subckt 1088_7443082010B_0.1u  1 2
Rp 1 2 29.46
Cp 1 2 46.22p
Rs 1 N3 0.000114
L1 N3 2 0.109u
.ends 1088_7443082010B_0.1u 
*******
.subckt 1088_7443082012_0.12u  1 2
Rp 1 2 38.47
Cp 1 2 40.99p
Rs 1 N3 0.00018
L1 N3 2 0.11975u
.ends 1088_7443082012_0.12u 
*******
.subckt 1088_7443082012B_0.12u  1 2
Rp 1 2 30.59
Cp 1 2 55.52p
Rs 1 N3 0.000114
L1 N3 2 0.128u
.ends 1088_7443082012B_0.12u 
*******
.subckt 1088_7443082015_0.15u  1 2
Rp 1 2 31.74
Cp 1 2 45.52p
Rs 1 N3 0.00018
L1 N3 2 0.13987u
.ends 1088_7443082015_0.15u 
*******
.subckt 1088_7443082015A_0.15u  1 2
Rp 1 2 33.62
Cp 1 2 54.7p
Rs 1 N3 0.00015
L1 N3 2 0.14707u
.ends 1088_7443082015A_0.15u 
*******
.subckt 1088_7443082015B_0.15u  1 2
Rp 1 2 32.09
Cp 1 2 62.84p
Rs 1 N3 0.000114
L1 N3 2 0.161u
.ends 1088_7443082015B_0.15u 
*******
.subckt 1088_7443082017_0.17u  1 2
Rp 1 2 30
Cp 1 2 57.6p
Rs 1 N3 0.00018
L1 N3 2 0.17644u
.ends 1088_7443082017_0.17u 
*******
.subckt 1088_7443082018_0.18u  1 2
Rp 1 2 30.33
Cp 1 2 44.82p
Rs 1 N3 0.00018
L1 N3 2 0.1795u
.ends 1088_7443082018_0.18u 
*******
.subckt 1088_7443082018A_0.18u  1 2
Rp 1 2 36.81
Cp 1 2 63.02p
Rs 1 N3 0.00015
L1 N3 2 0.18133u
.ends 1088_7443082018A_0.18u 
*******
.subckt 1088_7443082022_0.22u  1 2
Rp 1 2 33.66
Cp 1 2 53.18p
Rs 1 N3 0.00018
L1 N3 2 0.21486u
.ends 1088_7443082022_0.22u 
*******
.subckt 1323_74431323012_0.12u  1 2
Rp 1 2 67.84
Cp 1 2 3.53p
Rs 1 N3 0.00076
L1 N3 2 0.11974u
.ends 1323_74431323012_0.12u 
*******
.subckt 1323_74431323016_0.16u  1 2
Rp 1 2 66.58
Cp 1 2 10.29p
Rs 1 N3 0.00076
L1 N3 2 0.16128u
.ends 1323_74431323016_0.16u 
*******
.subckt 1411_7443091062_0.62u  1 2
Rp 1 2 59
Cp 1 2 69p
Rs 1 N3 0.00042
L1 N3 2 0.598u
.ends 1411_7443091062_0.62u 
*******
.subckt 1411_7443091080_0.8u  1 2
Rp 1 2 79
Cp 1 2 96p
Rs 1 N3 0.00042
L1 N3 2 0.767u
.ends 1411_7443091080_0.8u 
*******
.subckt 1411_7443091100_1u  1 2
Rp 1 2 103
Cp 1 2 57p
Rs 1 N3 0.00042
L1 N3 2 1u
.ends 1411_7443091100_1u 
*******
.subckt 1411_7443091120_1.2u  1 2
Rp 1 2 104
Cp 1 2 104p
Rs 1 N3 0.00042
L1 N3 2 1.2u
.ends 1411_7443091120_1.2u 
*******
.subckt 1411_7443091150_1.5u  1 2
Rp 1 2 107
Cp 1 2 93p
Rs 1 N3 0.00042
L1 N3 2 1.5u
.ends 1411_7443091150_1.5u 
*******
.subckt 1435_74431435010_0.1u  1 2
Rp 1 2 48
Cp 1 2 99p
Rs 1 N3 0.00028
L1 N3 2 0.106u
.ends 1435_74431435010_0.1u 
*******
.subckt 1435_74431435012_0.12u  1 2
Rp 1 2 51
Cp 1 2 134.6p
Rs 1 N3 0.00028
L1 N3 2 0.134u
.ends 1435_74431435012_0.12u 
*******
.subckt 1435_74431435015_0.15u  1 2
Rp 1 2 46
Cp 1 2 23p
Rs 1 N3 0.00028
L1 N3 2 0.148u
.ends 1435_74431435015_0.15u 
*******
.subckt 1435_74431435018_0.18u  1 2
Rp 1 2 52
Cp 1 2 32p
Rs 1 N3 0.00028
L1 N3 2 0.198u
.ends 1435_74431435018_0.18u 
*******
.subckt 1435_74431435022_0.22u  1 2
Rp 1 2 52
Cp 1 2 32p
Rs 1 N3 0.00028
L1 N3 2 0.224u
.ends 1435_74431435022_0.22u 
*******
.subckt 1435_74431435047_470n  1 2
Rp 1 2 54.433
Cp 1 2 50.806p
Rs 1 N3 0.00028
L1 N3 2 0.51001u
.ends 1435_74431435047_470n 
*******
.subckt 1012_74431012007_70n  1 2
Rp 1 2 41.444
Cp 1 2 7.467p
Rs 1 N3 0.000125
L1 N3 2 0.074731u
.ends 1012_74431012007_70n 
*******
.subckt 1012_74431012010_100n  1 2
Rp 1 2 33.974
Cp 1 2 35.541p
Rs 1 N3 0.000125
L1 N3 2 0.099838u
.ends 1012_74431012010_100n 
*******
.subckt 1012_74431012012_120n  1 2
Rp 1 2 37.049
Cp 1 2 34.381p
Rs 1 N3 0.000125
L1 N3 2 0.130404u
.ends 1012_74431012012_120n 
*******
.subckt 1012_74431012015_150n  1 2
Rp 1 2 41.646
Cp 1 2 33.261p
Rs 1 N3 0.000125
L1 N3 2 0.151517u
.ends 1012_74431012015_150n 
*******
.subckt 4030_744340300025_25n  1 2
Rp 1 2 23.5
Cp 1 2 24p
Rs 1 N3 0.0003105
L1 N3 2 0.025u
.ends 4030_744340300025_25n 
*******
.subckt 4030_744340300055_55n  1 2
Rp 1 2 29.321
Cp 1 2 29.299p
Rs 1 N3 0.0003105
L1 N3 2 0.056324u
.ends 4030_744340300055_55n 
*******
.subckt 4030_744340300075_75n  1 2
Rp 1 2 31.127
Cp 1 2 34.644p
Rs 1 N3 0.0003105
L1 N3 2 0.064746u
.ends 4030_744340300075_75n 
*******
.subckt 4035_74434035010_100n  1 2
Rp 1 2 31.361
Cp 1 2 58.945p
Rs 1 N3 0.00031
L1 N3 2 0.08684u
.ends 4035_74434035010_100n 
*******
.subckt 5030_74435030010_100n  1 2
Rp 1 2 37.557
Cp 1 2 37.678p
Rs 1 N3 0.0003565
L1 N3 2 0.096909u
.ends 5030_74435030010_100n 
*******
.subckt 9065_744300006_60n  1 2
Rp 1 2 27.774
Cp 1 2 26.65p
Rs 1 N3 0.00055
L1 N3 2 0.061889u
.ends 9065_744300006_60n 
*******
.subckt 9065_744300008_80n  1 2
Rp 1 2 28.724
Cp 1 2 36.05p
Rs 1 N3 0.00055
L1 N3 2 0.078758u
.ends 9065_744300008_80n 
*******
.subckt 9065_744300010_100n  1 2
Rp 1 2 30.193
Cp 1 2 46.623p
Rs 1 N3 0.00055
L1 N3 2 0.098291u
.ends 9065_744300010_100n 
*******
.subckt 9065_744300015_150n  1 2
Rp 1 2 33.62
Cp 1 2 67.437p
Rs 1 N3 0.002
L1 N3 2 0.146178u
.ends 9065_744300015_150n 
*******
.subckt 9065_744300022_220n  1 2
Rp 1 2 34.612
Cp 1 2 80.172p
Rs 1 N3 0.00055
L1 N3 2 0.218406u
.ends 9065_744300022_220n 
*******
.subckt 4035_74434035007_70n  1 2
Rp 1 2 26.7
Cp 1 2 51.328p
Rs 1 N3 0.00005
L1 N3 2 0.069035u
.ends 4035_74434035007_70n 
*******
.subckt 4030_744340300030_30n  1 2
Rp 1 2 21
Cp 1 2 25.328p
Rs 1 N3 0.085
L1 N3 2 0.023535u
.ends 4030_744340300030_30n 
*******
