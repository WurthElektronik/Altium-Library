**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ATUL
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 860040272001_100uF 1 2
Rser 1 3 0.20517788295
Lser 2 4 4.549671789E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860040272001_100uF
*******
.subckt 860040273002_220uF 1 2
Rser 1 3 0.12
Lser 2 4 0.0000000025
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860040273002_220uF
*******
.subckt 860040273003_330uF 1 2
Rser 1 3 0.09864
Lser 2 4 8.945178032E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860040273003_330uF
*******
.subckt 860040274004_470uF 1 2
Rser 1 3 0.068
Lser 2 4 0.000000007
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040274004_470uF
*******
.subckt 860040274005_680uF 1 2
Rser 1 3 0.05
Lser 2 4 0.000000011
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860040274005_680uF
*******
.subckt 860040274008_1mF 1 2
Rser 1 3 0.036
Lser 2 4 0.0000000025
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040274008_1mF
*******
.subckt 860040275006_680uF 1 2
Rser 1 3 0.042
Lser 2 4 0.000000007
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860040275006_680uF
*******
.subckt 860040275007_820uF 1 2
Rser 1 3 0.0345070171849
Lser 2 4 6.852542219E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860040275007_820uF
*******
.subckt 860040275009_1mF 1 2
Rser 1 3 0.034
Lser 2 4 0.000000006
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040275009_1mF
*******
.subckt 860040275010_1.2mF 1 2
Rser 1 3 0.0255844129341
Lser 2 4 9.696368316E-09
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860040275010_1.2mF
*******
.subckt 860040275011_1.5mF 1 2
Rser 1 3 0.022044936113
Lser 2 4 6.948768619E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860040275011_1.5mF
*******
.subckt 860040275012_2.2mF 1 2
Rser 1 3 0.0157262224146
Lser 2 4 5.66542288E-09
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860040275012_2.2mF
*******
.subckt 860040278013_2.2mF 1 2
Rser 1 3 0.022216481395
Lser 2 4 7.459394709E-09
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860040278013_2.2mF
*******
.subckt 860040278014_3.3mF 1 2
Rser 1 3 0.0212678160824
Lser 2 4 1.0398507261E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860040278014_3.3mF
*******
.subckt 860040278015_3.9mF 1 2
Rser 1 3 0.0164162128342
Lser 2 4 1.0766822979E-08
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860040278015_3.9mF
*******
.subckt 860040372001_56uF 1 2
Rser 1 3 0.2
Lser 2 4 0.000000002
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860040372001_56uF
*******
.subckt 860040373002_100uF 1 2
Rser 1 3 0.11
Lser 2 4 0.0000000035
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860040373002_100uF
*******
.subckt 860040373003_120uF 1 2
Rser 1 3 0.1
Lser 2 4 0.000000004
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860040373003_120uF
*******
.subckt 860040374004_220uF 1 2
Rser 1 3 0.08
Lser 2 4 0.000000004
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860040374004_220uF
*******
.subckt 860040374005_330uF 1 2
Rser 1 3 0.055
Lser 2 4 0.000000006
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860040374005_330uF
*******
.subckt 860040374006_470uF 1 2
Rser 1 3 0.0391400434095
Lser 2 4 5.417592351E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040374006_470uF
*******
.subckt 860040374008_680uF 1 2
Rser 1 3 0.039
Lser 2 4 0.000000004
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860040374008_680uF
*******
.subckt 860040375007_470uF 1 2
Rser 1 3 0.047
Lser 2 4 0.000000006
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040375007_470uF
*******
.subckt 860040375009_820uF 1 2
Rser 1 3 0.026
Lser 2 4 6.89756253077295E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860040375009_820uF
*******
.subckt 860040375010_1mF 1 2
Rser 1 3 0.0231016082725
Lser 2 4 7.51340742E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040375010_1mF
*******
.subckt 860040375012_1.2mF 1 2
Rser 1 3 0.0188603888594
Lser 2 4 7.418284491E-09
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860040375012_1.2mF
*******
.subckt 860040378011_1mF 1 2
Rser 1 3 0.0287553379109
Lser 2 4 9.175755509E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040378011_1mF
*******
.subckt 860040378013_1.5mF 1 2
Rser 1 3 0.0189631309012
Lser 2 4 6.875169541E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860040378013_1.5mF
*******
.subckt 860040378014_1.8mF 1 2
Rser 1 3 0.0174527376895
Lser 2 4 9.271190652E-09
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860040378014_1.8mF
*******
.subckt 860040378015_2.2mF 1 2
Rser 1 3 0.0197044613681
Lser 2 4 8.826746349E-09
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860040378015_2.2mF
*******
.subckt 860040378016_2.7mF 1 2
Rser 1 3 0.0150102484108
Lser 2 4 8.489873224E-09
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860040378016_2.7mF
*******
.subckt 860040378017_3.3mF 1 2
Rser 1 3 0.014212785855
Lser 2 4 1.0973141819E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860040378017_3.3mF
*******
.subckt 860040381018_4.7mF 1 2
Rser 1 3 0.0169941417717
Lser 2 4 1.9483441233E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860040381018_4.7mF
*******
.subckt 860040472001_47uF 1 2
Rser 1 3 0.236760667715
Lser 2 4 5.219330547E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860040472001_47uF
*******
.subckt 860040472002_56uF 1 2
Rser 1 3 0.148
Lser 2 4 0.0000000025
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860040472002_56uF
*******
.subckt 860040473003_100uF 1 2
Rser 1 3 0.0909990443008
Lser 2 4 3.859469302E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860040473003_100uF
*******
.subckt 860040474004_220uF 1 2
Rser 1 3 0.08
Lser 2 4 0.000000023
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860040474004_220uF
*******
.subckt 860040474005_330uF 1 2
Rser 1 3 0.048
Lser 2 4 0.000000011
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860040474005_330uF
*******
.subckt 860040474007_470uF 1 2
Rser 1 3 0.033
Lser 2 4 0.000000009
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040474007_470uF
*******
.subckt 860040475006_330uF 1 2
Rser 1 3 0.044
Lser 2 4 0.000000004
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860040475006_330uF
*******
.subckt 860040475008_470uF 1 2
Rser 1 3 0.035
Lser 2 4 0.000000008
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040475008_470uF
*******
.subckt 860040475009_680uF 1 2
Rser 1 3 0.0230221005822
Lser 2 4 5.921120681E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860040475009_680uF
*******
.subckt 860040475010_820uF 1 2
Rser 1 3 0.0190009846867
Lser 2 4 5.849771069E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860040475010_820uF
*******
.subckt 860040475011_1mF 1 2
Rser 1 3 0.0205234255636
Lser 2 4 6.33869368E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040475011_1mF
*******
.subckt 860040478012_1mF 1 2
Rser 1 3 0.0208810202664
Lser 2 4 6.126211991E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040478012_1mF
*******
.subckt 860040478013_1.5mF 1 2
Rser 1 3 0.0180672352148
Lser 2 4 9.793779097E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860040478013_1.5mF
*******
.subckt 860040478014_1.8mF 1 2
Rser 1 3 0.0163859824822
Lser 2 4 8.815281386E-09
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860040478014_1.8mF
*******
.subckt 860040478015_2.2mF 1 2
Rser 1 3 0.0117488115195
Lser 2 4 9.492955498E-09
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860040478015_2.2mF
*******
.subckt 860040480016_2.7mF 1 2
Rser 1 3 0.0175427236178
Lser 2 4 1.7730717395E-08
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860040480016_2.7mF
*******
.subckt 860040572001_33uF 1 2
Rser 1 3 0.19
Lser 2 4 0.000000003
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860040572001_33uF
*******
.subckt 860040572002_47uF 1 2
Rser 1 3 0.175
Lser 2 4 0.000000002
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860040572002_47uF
*******
.subckt 860040573003_56uF 1 2
Rser 1 3 0.127
Lser 2 4 0.0000000045
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860040573003_56uF
*******
.subckt 860040573004_100uF 1 2
Rser 1 3 0.1
Lser 2 4 0.0000000035
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860040573004_100uF
*******
.subckt 860040574005_150uF 1 2
Rser 1 3 0.068
Lser 2 4 0.000000009
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860040574005_150uF
*******
.subckt 860040574006_220uF 1 2
Rser 1 3 0.0483035818626
Lser 2 4 4.633219958E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860040574006_220uF
*******
.subckt 860040574008_270uF 1 2
Rser 1 3 0.038
Lser 2 4 0.000000005
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860040574008_270uF
*******
.subckt 860040575007_220uF 1 2
Rser 1 3 0.052
Lser 2 4 0.000000009
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860040575007_220uF
*******
.subckt 860040575009_330uF 1 2
Rser 1 3 0.037
Lser 2 4 0.000000011
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860040575009_330uF
*******
.subckt 860040575010_470uF 1 2
Rser 1 3 0.0231728091811
Lser 2 4 7.713499455E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040575010_470uF
*******
.subckt 860040575011_560uF 1 2
Rser 1 3 0.0211825859338
Lser 2 4 5.875444861E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860040575011_560uF
*******
.subckt 860040575012_680uF 1 2
Rser 1 3 0.0183533764035
Lser 2 4 7.462454355E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860040575012_680uF
*******
.subckt 860040578013_680uF 1 2
Rser 1 3 0.0235127310626
Lser 2 4 8.946424739E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860040578013_680uF
*******
.subckt 860040578014_1mF 1 2
Rser 1 3 0.020010707593
Lser 2 4 8.222422508E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040578014_1mF
*******
.subckt 860040578015_1.2mF 1 2
Rser 1 3 0.0163465169374
Lser 2 4 8.811463148E-09
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860040578015_1.2mF
*******
.subckt 860040578017_1.5mF 1 2
Rser 1 3 0.0133840092478
Lser 2 4 9.396241494E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860040578017_1.5mF
*******
.subckt 860040580016_1.2mF 1 2
Rser 1 3 0.018966462855
Lser 2 4 1.7114535337E-08
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860040580016_1.2mF
*******
.subckt 860040580018_1.8mF 1 2
Rser 1 3 0.0198457933443
Lser 2 4 1.4245271502E-08
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860040580018_1.8mF
*******
.subckt 860040580019_2.7mF 1 2
Rser 1 3 0.0127605149046
Lser 2 4 1.5725414079E-08
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860040580019_2.7mF
*******
.subckt 860040581020_2.7mF 1 2
Rser 1 3 0.0166495852009
Lser 2 4 1.7201267115E-08
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860040581020_2.7mF
*******
.subckt 860040581021_4.7mF 1 2
Rser 1 3 0.015
Lser 2 4 0.00000001
C1 3 4 0.0047
Rpar 3 4 21276.5957446808
.ends 860040581021_4.7mF
*******
.subckt 860040672001_22uF 1 2
Rser 1 3 0.23
Lser 2 4 0.000000003
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860040672001_22uF
*******
.subckt 860040673002_47uF 1 2
Rser 1 3 0.25
Lser 2 4 0.000000003
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860040673002_47uF
*******
.subckt 860040673003_56uF 1 2
Rser 1 3 0.087
Lser 2 4 0.000000006
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860040673003_56uF
*******
.subckt 860040674004_100uF 1 2
Rser 1 3 0.1
Lser 2 4 0.0000000205
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860040674004_100uF
*******
.subckt 860040674005_120uF 1 2
Rser 1 3 0.058
Lser 2 4 0.000000008
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860040674005_120uF
*******
.subckt 860040674007_180uF 1 2
Rser 1 3 0.046
Lser 2 4 0.000000006
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860040674007_180uF
*******
.subckt 860040675006_150uF 1 2
Rser 1 3 0.0489086457007
Lser 2 4 6.882764417E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860040675006_150uF
*******
.subckt 860040675008_220uF 1 2
Rser 1 3 0.042
Lser 2 4 0.00000001
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860040675008_220uF
*******
.subckt 860040675009_270uF 1 2
Rser 1 3 0.0270499784263
Lser 2 4 7.797139219E-09
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860040675009_270uF
*******
.subckt 860040675010_330uF 1 2
Rser 1 3 0.0236848215901
Lser 2 4 5.647450413E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860040675010_330uF
*******
.subckt 860040675011_470uF 1 2
Rser 1 3 0.045
Lser 2 4 0.000000007
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040675011_470uF
*******
.subckt 860040678012_560uF 1 2
Rser 1 3 0.0197171314895
Lser 2 4 7.858123212E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860040678012_560uF
*******
.subckt 860040680013_1.2mF 1 2
Rser 1 3 0.0366474562282
Lser 2 4 1.5684772409E-08
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860040680013_1.2mF
*******
.subckt 860040773001_33uF 1 2
Rser 1 3 0.578633024315
Lser 2 4 4.618903108E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860040773001_33uF
*******
.subckt 860040774002_47uF 1 2
Rser 1 3 0.18
Lser 2 4 0.0000000045
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860040774002_47uF
*******
.subckt 860040774003_56uF 1 2
Rser 1 3 0.15
Lser 2 4 0.000000006
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860040774003_56uF
*******
.subckt 860040774004_82uF 1 2
Rser 1 3 0.165
Lser 2 4 0.0000000045
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860040774004_82uF
*******
.subckt 860040774007_120uF 1 2
Rser 1 3 0.13
Lser 2 4 0.000000004
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860040774007_120uF
*******
.subckt 860040775005_82uF 1 2
Rser 1 3 0.154
Lser 2 4 0.000000005
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860040775005_82uF
*******
.subckt 860040775006_100uF 1 2
Rser 1 3 0.18
Lser 2 4 0.0000000035
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860040775006_100uF
*******
.subckt 860040775008_120uF 1 2
Rser 1 3 0.105
Lser 2 4 0.000000008
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860040775008_120uF
*******
.subckt 860040775009_180uF 1 2
Rser 1 3 0.107
Lser 2 4 0.000000005
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860040775009_180uF
*******
.subckt 860040775010_220uF 1 2
Rser 1 3 0.048
Lser 2 4 0.000000007
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860040775010_220uF
*******
.subckt 860040778011_270uF 1 2
Rser 1 3 0.0729917824506
Lser 2 4 7.997228003E-09
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860040778011_270uF
*******
.subckt 860040778012_330uF 1 2
Rser 1 3 0.064
Lser 2 4 0.000000011
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860040778012_330uF
*******
.subckt 860040778013_470uF 1 2
Rser 1 3 0.055
Lser 2 4 0.000000013
C1 3 4 0.00047
Rpar 3 4 212765.957446808
.ends 860040778013_470uF
*******
.subckt 860040778015_680uF 1 2
Rser 1 3 0.041
Lser 2 4 0.00000003
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860040778015_680uF
*******
.subckt 860040780014_560uF 1 2
Rser 1 3 0.048
Lser 2 4 0.000000007
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860040780014_560uF
*******
.subckt 860040780016_820uF 1 2
Rser 1 3 0.0225
Lser 2 4 0.000000015
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860040780016_820uF
*******
.subckt 860040780017_1mF 1 2
Rser 1 3 0.0296677915498
Lser 2 4 1.6402235434E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040780017_1mF
*******
.subckt 860040780019_1.2mF 1 2
Rser 1 3 0.034
Lser 2 4 0.000000028
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860040780019_1.2mF
*******
.subckt 860040781018_1mF 1 2
Rser 1 3 0.0312938724538
Lser 2 4 1.3804216007E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 860040781018_1mF
*******
.subckt 860040781020_1.2mF 1 2
Rser 1 3 0.023671459975
Lser 2 4 1.6482381522E-08
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860040781020_1.2mF
*******
.subckt 860040781021_1.5mF 1 2
Rser 1 3 0.0242402948837
Lser 2 4 1.6980212185E-08
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860040781021_1.5mF
*******
.subckt 860040874001_27uF 1 2
Rser 1 3 0.416549391839
Lser 2 4 4.070972199E-09
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 860040874001_27uF
*******
.subckt 860040875002_47uF 1 2
Rser 1 3 0.234056685461
Lser 2 4 5.361797892E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860040875002_47uF
*******
.subckt 860040875003_68uF 1 2
Rser 1 3 0.152
Lser 2 4 0.000000004
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860040875003_68uF
*******
.subckt 860040875004_82uF 1 2
Rser 1 3 0.073
Lser 2 4 0.000000009
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860040875004_82uF
*******
.subckt 860040875005_100uF 1 2
Rser 1 3 0.144
Lser 2 4 0.000000005
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860040875005_100uF
*******
.subckt 860040878006_120uF 1 2
Rser 1 3 0.0768083693712
Lser 2 4 6.761056573E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860040878006_120uF
*******
.subckt 860040878008_330uF 1 2
Rser 1 3 0.0301199755611
Lser 2 4 8.796266061E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860040878008_330uF
*******
.subckt 860040880007_270uF 1 2
Rser 1 3 0.052
Lser 2 4 0.000000011
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860040880007_270uF
*******
.subckt 860040880009_390uF 1 2
Rser 1 3 0.039748091695
Lser 2 4 1.57277015E-08
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860040880009_390uF
*******
.subckt 860040880011_470uF 1 2
Rser 1 3 0.036
Lser 2 4 0.000000011
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040880011_470uF
*******
.subckt 860040881010_390uF 1 2
Rser 1 3 0.0472471077084
Lser 2 4 1.6544964659E-08
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860040881010_390uF
*******
.subckt 860040881012_470uF 1 2
Rser 1 3 0.04
Lser 2 4 0.000000009
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860040881012_470uF
*******
.subckt 860040881013_680uF 1 2
Rser 1 3 0.0312965081231
Lser 2 4 1.4954980575E-08
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860040881013_680uF
*******
.subckt 860040881014_820uF 1 2
Rser 1 3 0.0296245810975
Lser 2 4 1.4842917536E-08
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860040881014_820uF
*******
