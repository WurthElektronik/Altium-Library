**************************************************
* Manufacturer:          Würth Elektronik
* Kinds:                 SMT Shielded Power Inductor
* Matchcode:             WE-PDA
* Library Type:          LTspice
* Version:               rev23a
* Created/modified by:   Ella
* Date and Time:         8/7/2023
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2023 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 1210_7847709010_1u 1 2
Rp 1 2 2294.915406849
Cp 1 2 1.3882750261p
Rs 1 N3 0.008
L1 N3 2 0.9477912049945u
.ends 1210_7847709010_1u
*******
.subckt 1210_7847709022_2.2u 1 2
Rp 1 2 4769.985971776
Cp 1 2 1.5093643078p
Rs 1 N3 0.012
L1 N3 2 2.265509355663u
.ends 1210_7847709022_2.2u
*******
.subckt 1210_7847709033_3.3u 1 2
Rp 1 2 6338.363617445
Cp 1 2 1.6117205723p
Rs 1 N3 0.014
L1 N3 2 3.116581080998u
.ends 1210_7847709033_3.3u
*******
.subckt 1210_7847709047_4.7u 1 2
Rp 1 2 7853.568425335
Cp 1 2 1.7532943876p
Rs 1 N3 0.016
L1 N3 2 4.11518615215u
.ends 1210_7847709047_4.7u
*******
.subckt 1210_7847709068_6.8u 1 2
Rp 1 2 11244.49787969
Cp 1 2 2.7755980227p
Rs 1 N3 0.02
L1 N3 2 6.380294136413u
.ends 1210_7847709068_6.8u
*******
.subckt 1210_7847709100_10u 1 2
Rp 1 2 14651.33471798
Cp 1 2 5.1433007426p
Rs 1 N3 0.025
L1 N3 2 9.454216640987u
.ends 1210_7847709100_10u
*******
.subckt 1210_7847709150_15u 1 2
Rp 1 2 19799
Cp 1 2 3.95p
Rs 1 N3 0.03
L1 N3 2 14.93u
.ends 1210_7847709150_15u
*******
.subckt 1210_7847709220_22u 1 2
Rp 1 2 24529.7119385
Cp 1 2 9.1256019813p
Rs 1 N3 0.037
L1 N3 2 19.49383174863u
.ends 1210_7847709220_22u
*******
.subckt 1210_7847709330_33u 1 2
Rp 1 2 26829
Cp 1 2 10.3p
Rs 1 N3 0.0443
L1 N3 2 29.924u
.ends 1210_7847709330_33u
*******
.subckt 1210_7847709470_47u 1 2
Rp 1 2 46246.28473571
Cp 1 2 15.428751801p
Rs 1 N3 0.056
L1 N3 2 41.90253832625u
.ends 1210_7847709470_47u
*******
.subckt 1210_7847709680_68u 1 2
Rp 1 2 59363
Cp 1 2 11.8p
Rs 1 N3 0.0655
L1 N3 2 62.137u
.ends 1210_7847709680_68u
*******
.subckt 1210_7847709101_100u 1 2
Rp 1 2 101541.0668698
Cp 1 2 12.7073566505p
Rs 1 N3 0.1
L1 N3 2 87.16698574827u
.ends 1210_7847709101_100u
*******
.subckt 1210_7847709221_220u 1 2
Rp 1 2 105097.46965648
Cp 1 2 16.0315674238p
Rs 1 N3 0.205
L1 N3 2 196.7291808281u
.ends 1210_7847709221_220u
*******
.subckt 1210_7847709331_330u 1 2
Rp 1 2 89155
Cp 1 2 17p
Rs 1 N3 0.34
L1 N3 2 319.916u
.ends 1210_7847709331_330u
*******
.subckt 1210_7847709471_470u 1 2
Rp 1 2 109394.88869077
Cp 1 2 17.578119258p
Rs 1 N3 0.41
L1 N3 2 390.1587144886u
.ends 1210_7847709471_470u
*******
.subckt 1210_7847709102_1000u 1 2
Rp 1 2 216540.591668429
Cp 1 2 15.7632287615714p
Rs 1 N3 0.885
L1 N3 2 774.510514956553u
.ends 1210_7847709102_1000u
*******
.subckt 1260_784771010_1u 1 2
Rp 1 2 2433.248526684
Cp 1 2 1.3484119846p
Rs 1 N3 0.007
L1 N3 2 0.964037u
.ends 1260_784771010_1u
*******
.subckt 1260_784771022_2.2u 1 2
Rp 1 2 5189.569854217
Cp 1 2 1.6159803997p
Rs 1 N3 0.0105
L1 N3 2 2.292796219119u
.ends 1260_784771022_2.2u
*******
.subckt 1260_784771033_3.3u 1 2
Rp 1 2 7131.108427517
Cp 1 2 1.6514667945p
Rs 1 N3 0.012
L1 N3 2 3.24701584243u
.ends 1260_784771033_3.3u
*******
.subckt 1260_784771047_4.7u 1 2
Rp 1 2 9042.156448366
Cp 1 2 2.4368902869p
Rs 1 N3 0.0145
L1 N3 2 4.261980332565u
.ends 1260_784771047_4.7u
*******
.subckt 1260_784771068_6.8u 1 2
Rp 1 2 12513.50740286
Cp 1 2 4.8563450773p
Rs 1 N3 0.018
L1 N3 2 6.824458759468u
.ends 1260_784771068_6.8u
*******
.subckt 1260_784771082_8.2u 1 2
Rp 1 2 14787.17407293
Cp 1 2 4.8158190373p
Rs 1 N3 0.02
L1 N3 2 8.274635790997u
.ends 1260_784771082_8.2u
*******
.subckt 1260_784771100_10u 1 2
Rp 1 2 17178.30402294
Cp 1 2 5.2969598266p
Rs 1 N3 0.022
L1 N3 2 9.854886153843u
.ends 1260_784771100_10u
*******
.subckt 1260_784771220_22u 1 2
Rp 1 2 31803.37051151
Cp 1 2 5.8357084029p
Rs 1 N3 0.0335
L1 N3 2 19.61866271393u
.ends 1260_784771220_22u
*******
.subckt 1260_784771330_33u 1 2
Rp 1 2 40694
Cp 1 2 6.2p
Rs 1 N3 0.052
L1 N3 2 30.717u
.ends 1260_784771330_33u
*******
.subckt 1260_784771470_47u 1 2
Rp 1 2 52452.11268997
Cp 1 2 6.1761314516p
Rs 1 N3 0.064
L1 N3 2 40.5429765455u
.ends 1260_784771470_47u
*******
.subckt 1260_784771680_68u 1 2
Rp 1 2 65310
Cp 1 2 5.9p
Rs 1 N3 0.115
L1 N3 2 65.472u
.ends 1260_784771680_68u
*******
.subckt 1260_784771101_100u 1 2
Rp 1 2 96751.83862672
Cp 1 2 6.6698797519p
Rs 1 N3 0.145
L1 N3 2 89.45051933212u
.ends 1260_784771101_100u
*******
.subckt 1260_784771221_220u 1 2
Rp 1 2 105001.69441514
Cp 1 2 8.886001314p
Rs 1 N3 0.29
L1 N3 2 189.7638052611u
.ends 1260_784771221_220u
*******
.subckt 1260_784771331_330u 1 2
Rp 1 2 254752
Cp 1 2 7.56p
Rs 1 N3 0.495
L1 N3 2 314.264u
.ends 1260_784771331_330u
*******
.subckt 1260_784771471_470u 1 2
Rp 1 2 251375.1912763
Cp 1 2 6.5663338599p
Rs 1 N3 0.588
L1 N3 2 439.2246612792u
.ends 1260_784771471_470u
*******
.subckt 1260_784771102_1000u 1 2
Rp 1 2 184405.7372337
Cp 1 2 8.9931636428p
Rs 1 N3 1.42
L1 N3 2 958.0309208405u
.ends 1260_784771102_1000u
*******
.subckt 1280_78477010_1u 1 2
Rp 1 2 2668.882619536
Cp 1 2 1.2949025235p
Rs 1 N3 0.0075
L1 N3 2 0.851361u
.ends 1280_78477010_1u
*******
.subckt 1280_78477022_2.2u 1 2
Rp 1 2 5813.474815798
Cp 1 2 1.5220075628p
Rs 1 N3 0.012
L1 N3 2 2.286935796312u
.ends 1280_78477022_2.2u
*******
.subckt 1280_78477033_3.3u 1 2
Rp 1 2 7614.617238701
Cp 1 2 1.5416464406p
Rs 1 N3 0.014
L1 N3 2 3.212340743703u
.ends 1280_78477033_3.3u
*******
.subckt 1280_78477047_4.7u 1 2
Rp 1 2 9407.872771631
Cp 1 2 1.7999782823p
Rs 1 N3 0.0165
L1 N3 2 4.206935362839u
.ends 1280_78477047_4.7u
*******
.subckt 1280_78477068_6.8u 1 2
Rp 1 2 14556.74736043
Cp 1 2 2.1384636392p
Rs 1 N3 0.021
L1 N3 2 6.798057276949u
.ends 1280_78477068_6.8u
*******
.subckt 1280_784770100_10u 1 2
Rp 1 2 18808.39861138
Cp 1 2 3.2660671847p
Rs 1 N3 0.026
L1 N3 2 9.940123740059u
.ends 1280_784770100_10u
*******
.subckt 1280_784770220_22u 1 2
Rp 1 2 31940.81996524
Cp 1 2 5.2589619092p
Rs 1 N3 0.037
L1 N3 2 20.19197852179u
.ends 1280_784770220_22u
*******
.subckt 1280_784770330_33u 1 2
Rp 1 2 25921
Cp 1 2 9.75p
Rs 1 N3 0.0458
L1 N3 2 29.022u
.ends 1280_784770330_33u
*******
.subckt 1280_784770470_47u 1 2
Rp 1 2 56578.20721198
Cp 1 2 9.5024623536p
Rs 1 N3 0.059
L1 N3 2 42.7394983986u
.ends 1280_784770470_47u
*******
.subckt 1280_784770680_68u 1 2
Rp 1 2 72516
Cp 1 2 9.849p
Rs 1 N3 0.082
L1 N3 2 64.774u
.ends 1280_784770680_68u
*******
.subckt 1280_784770101_100u 1 2
Rp 1 2 97590.86624169
Cp 1 2 10.4463930828p
Rs 1 N3 0.12
L1 N3 2 92.07199101756u
.ends 1280_784770101_100u
*******
.subckt 1280_784770221_220u 1 2
Rp 1 2 133347.06902775
Cp 1 2 11.2068371226p
Rs 1 N3 0.25
L1 N3 2 207.6478051298u
.ends 1280_784770221_220u
*******
.subckt 1280_784770331_330u 1 2
Rp 1 2 364620
Cp 1 2 11.8p
Rs 1 N3 0.39
L1 N3 2 324.661u
.ends 1280_784770331_330u
*******
.subckt 1280_784770471_470u 1 2
Rp 1 2 145181.648050917
Cp 1 2 14.2376988305p
Rs 1 N3 0.475
L1 N3 2 426.004640068417u
.ends 1280_784770471_470u
*******
.subckt 1280_784770102_1000u 1 2
Rp 1 2 83224.4700293857
Cp 1 2 12.2029488045714p
Rs 1 N3 1
L1 N3 2 922.109905113286u
.ends 1280_784770102_1000u
*******
.subckt 7332_784778010_1u 1 2
Rp 1 2 2307.40930898667
Cp 1 2 0.911242807222222p
Rs 1 N3 0.03
L1 N3 2 0.832000064693222u
.ends 7332_784778010_1u
*******
.subckt 7332_784778022_2.2u 1 2
Rp 1 2 4386.408048314
Cp 1 2 1.1974692155p
Rs 1 N3 0.042
L1 N3 2 1.718141625726u
.ends 7332_784778022_2.2u
*******
.subckt 7332_784778033_3.3u 1 2
Rp 1 2 6872.321544054
Cp 1 2 1.6662349176p
Rs 1 N3 0.054
L1 N3 2 3.004108330661u
.ends 7332_784778033_3.3u
*******
.subckt 7332_784778047_4.7u 1 2
Rp 1 2 9766.275617278
Cp 1 2 2.0898529192p
Rs 1 N3 0.066
L1 N3 2 4.589667711701u
.ends 7332_784778047_4.7u
*******
.subckt 7332_784778068_6.8u 1 2
Rp 1 2 13715.85350611
Cp 1 2 2.3775454772p
Rs 1 N3 0.079
L1 N3 2 6.499001324887u
.ends 7332_784778068_6.8u
*******
.subckt 7332_784778082_8.2u 1 2
Rp 1 2 15327.46241456
Cp 1 2 2.5060305278p
Rs 1 N3 0.086
L1 N3 2 7.602082540708u
.ends 7332_784778082_8.2u
*******
.subckt 7332_784778100_10u 1 2
Rp 1 2 19048.09163139
Cp 1 2 2.3265136356p
Rs 1 N3 0.105
L1 N3 2 9.76308112938u
.ends 7332_784778100_10u
*******
.subckt 7332_784778220_22u 1 2
Rp 1 2 14695.937803447
Cp 1 2 3.8904200749p
Rs 1 N3 0.156
L1 N3 2 21.35398943466u
.ends 7332_784778220_22u
*******
.subckt 7332_784778470_47u 1 2
Rp 1 2 61264.0585634545
Cp 1 2 3.19500997990909p
Rs 1 N3 0.29
L1 N3 2 44.2552423483909u
.ends 7332_784778470_47u
*******
.subckt 7332_784778101_100u 1 2
Rp 1 2 101282.362281329
Cp 1 2 3.28573847857143p
Rs 1 N3 0.6
L1 N3 2 90.9322883183429u
.ends 7332_784778101_100u
*******
.subckt 7332_784778221_220u 1 2
Rp 1 2 159660.763658714
Cp 1 2 3.38695254571429p
Rs 1 N3 1.35
L1 N3 2 196.783905129857u
.ends 7332_784778221_220u
*******
.subckt 7332_784778471_470u 1 2
Rp 1 2 231349.867191571
Cp 1 2 3.56735840542857p
Rs 1 N3 2.74
L1 N3 2 431.598145631286u
.ends 7332_784778471_470u
*******
.subckt 7332_784778102_1000u 1 2
Rp 1 2 389989
Cp 1 2 3.7085p
Rs 1 N3 6
L1 N3 2 896.011u
.ends 7332_784778102_1000u
*******
.subckt 7345_784777010_1u 1 2
Rp 1 2 2090.81936509
Cp 1 2 0.843162657p
Rs 1 N3 0.032
L1 N3 2 0.7836534724718u
.ends 7345_784777010_1u
*******
.subckt 7345_784777022_2.2u 1 2
Rp 1 2 4971.390102369
Cp 1 2 1.2907595592p
Rs 1 N3 0.051
L1 N3 2 2.180016129345u
.ends 7345_784777022_2.2u
*******
.subckt 7345_784777033_3.3u 1 2
Rp 1 2 6194.42616025222
Cp 1 2 1.202188746p
Rs 1 N3 0.058
L1 N3 2 2.76853435648111u
.ends 7345_784777033_3.3u
*******
.subckt 7345_784777047_4.7u 1 2
Rp 1 2 8557.586509961
Cp 1 2 1.4744181502p
Rs 1 N3 0.07
L1 N3 2 4.187187927039u
.ends 7345_784777047_4.7u
*******
.subckt 7345_784777068_6.8u 1 2
Rp 1 2 11500.66279623
Cp 1 2 1.9096557529p
Rs 1 N3 0.083
L1 N3 2 5.967935344578u
.ends 7345_784777068_6.8u
*******
.subckt 7345_784777082_8.2u 1 2
Rp 1 2 14719.48288191
Cp 1 2 2.3741500394p
Rs 1 N3 0.0975
L1 N3 2 7.895868403929u
.ends 7345_784777082_8.2u
*******
.subckt 7345_784777100_10u 1 2
Rp 1 2 15520.93335219
Cp 1 2 2.6257437707p
Rs 1 N3 0.105
L1 N3 2 9.111060714667u
.ends 7345_784777100_10u
*******
.subckt 7345_784777220_22u 1 2
Rp 1 2 34713.49948107
Cp 1 2 3.5868691419p
Rs 1 N3 0.18
L1 N3 2 21.0156666716u
.ends 7345_784777220_22u
*******
.subckt 7345_784777470_47u 1 2
Rp 1 2 39241.3504016
Cp 1 2 5.7367557873p
Rs 1 N3 0.25
L1 N3 2 42.93535458839u
.ends 7345_784777470_47u
*******
.subckt 7345_784777101_100u 1 2
Rp 1 2 70704.55918037
Cp 1 2 5.1165584441p
Rs 1 N3 0.39
L1 N3 2 88.06383986551u
.ends 7345_784777101_100u
*******
.subckt 7345_784777221_220u 1 2
Rp 1 2 100867.0948967
Cp 1 2 6.9140589382p
Rs 1 N3 0.945
L1 N3 2 199.7427916773u
.ends 7345_784777221_220u
*******
.subckt 7345_784777331_330u 1 2
Rp 1 2 203468
Cp 1 2 4.3p
Rs 1 N3 1.56
L1 N3 2 308.206u
.ends 7345_784777331_330u
*******
.subckt 7345_784777471_470u 1 2
Rp 1 2 177769.9360378
Cp 1 2 6.7437216173p
Rs 1 N3 2.27
L1 N3 2 443.9123496208u
.ends 7345_784777471_470u
*******
.subckt 7345_784777102_1000u 1 2
Rp 1 2 241276.825991857
Cp 1 2 8.166242278p
Rs 1 N3 4.8
L1 N3 2 910.643699477u
.ends 7345_784777102_1000u
*******
.subckt 1050_7847714033_3.3u 1 2
Rp 1 2 2007
Cp 1 2 9.206p
Rs 1 N3 0.012
L1 N3 2 3.271u
.ends 1050_7847714033_3.3u
*******
.subckt 1050_7847714047_4.7u 1 2
Rp 1 2 3886
Cp 1 2 9.489p
Rs 1 N3 0.014
L1 N3 2 4.189u
.ends 1050_7847714047_4.7u
*******
.subckt 1050_7847714100_10u 1 2
Rp 1 2 7924
Cp 1 2 10.391p
Rs 1 N3 0.026
L1 N3 2 8.684u
.ends 1050_7847714100_10u
*******
.subckt 1050_7847714220_22u 1 2
Rp 1 2 16615
Cp 1 2 12.333p
Rs 1 N3 0.063
L1 N3 2 22.297u
.ends 1050_7847714220_22u
*******
.subckt 1050_7847714330_33u 1 2
Rp 1 2 21893
Cp 1 2 11.489p
Rs 1 N3 0.079
L1 N3 2 31.318u
.ends 1050_7847714330_33u
*******
.subckt 1050_7847714470_47u 1 2
Rp 1 2 23438
Cp 1 2 13.651p
Rs 1 N3 0.123
L1 N3 2 45.46u
.ends 1050_7847714470_47u
*******
.subckt 1050_7847714680_68u 1 2
Rp 1 2 29832
Cp 1 2 13.617p
Rs 1 N3 0.147
L1 N3 2 60.755u
.ends 1050_7847714680_68u
*******
.subckt 1050_7847714101_100u 1 2
Rp 1 2 32869
Cp 1 2 14.482p
Rs 1 N3 0.245
L1 N3 2 90.064u
.ends 1050_7847714101_100u
*******
.subckt 1050_7847714221_220u 1 2
Rp 1 2 53359
Cp 1 2 14.021p
Rs 1 N3 0.59
L1 N3 2 214.773u
.ends 1050_7847714221_220u
*******
.subckt 1050_7847714331_330u 1 2
Rp 1 2 67719
Cp 1 2 13.604p
Rs 1 N3 0.75
L1 N3 2 318.302u
.ends 1050_7847714331_330u
*******
