**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Polymer Capacitors
* Matchcode:             WCAP-PSLC
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 875075155001_180uF 1 2
Rser 1 3 0.0135478480891
Lser 2 4 4.02110962E-09
C1 3 4 0.00018
Rpar 3 4 27777.7777777778
.ends 875075155001_180uF
*******
.subckt 875075155002_220uF 1 2
Rser 1 3 0.0062
Lser 2 4 0.000000004
C1 3 4 0.00022
Rpar 3 4 22727.2727272727
.ends 875075155002_220uF
*******
.subckt 875075155003_270uF 1 2
Rser 1 3 0.00499962712265
Lser 2 4 4.284889243E-09
C1 3 4 0.00027
Rpar 3 4 18518.5185185185
.ends 875075155003_270uF
*******
.subckt 875075155004_330uF 1 2
Rser 1 3 0.0064084536534
Lser 2 4 5.866294544E-09
C1 3 4 0.00033
Rpar 3 4 15144.2307692308
.ends 875075155004_330uF
*******
.subckt 875075155005_390uF 1 2
Rser 1 3 0.00518549626992
Lser 2 4 4.102648333E-09
C1 3 4 0.00039
Rpar 3 4 12830.9572301426
.ends 875075155005_390uF
*******
.subckt 875075155006_470uF 1 2
Rser 1 3 0.0073
Lser 2 4 0.0000000023
C1 3 4 0.00047
Rpar 3 4 10641.8918918919
.ends 875075155006_470uF
*******
.subckt 875075155008_680uF 1 2
Rser 1 3 0.00523627827166
Lser 2 4 4.046346351E-09
C1 3 4 0.00068
Rpar 3 4 7359.81308411215
.ends 875075155008_680uF
*******
.subckt 875075155009_820uF 1 2
Rser 1 3 0.00509349861377
Lser 2 4 3.981534221E-09
C1 3 4 0.00082
Rpar 3 4 6097.56097560976
.ends 875075155009_820uF
*******
.subckt 875075155010_1mF 1 2
Rser 1 3 0.00626328739571
Lser 2 4 4.179160925E-09
C1 3 4 0.001
Rpar 3 4 5000
.ends 875075155010_1mF
*******
.subckt 875075161011_1.2mF 1 2
Rser 1 3 0.00649673829676
Lser 2 4 5.37864984E-09
C1 3 4 0.0012
Rpar 3 4 4166.66666666667
.ends 875075161011_1.2mF
*******
.subckt 875075161012_1.5mF 1 2
Rser 1 3 0.00640729145682
Lser 2 4 5.168483696E-09
C1 3 4 0.0015
Rpar 3 4 3333.33333333333
.ends 875075161012_1.5mF
*******
.subckt 875075161013_2mF 1 2
Rser 1 3 0.0068215381043
Lser 2 4 5.301915109E-09
C1 3 4 0.002
Rpar 3 4 2500
.ends 875075161013_2mF
*******
.subckt 875075355001_180uF 1 2
Rser 1 3 0.0104669984726
Lser 2 4 3.95005494E-09
C1 3 4 0.00018
Rpar 3 4 27777.7777777778
.ends 875075355001_180uF
*******
.subckt 875075355002_220uF 1 2
Rser 1 3 0.0089594133143
Lser 2 4 3.977814839E-09
C1 3 4 0.00022
Rpar 3 4 22727.2727272727
.ends 875075355002_220uF
*******
.subckt 875075355003_270uF 1 2
Rser 1 3 0.00693451605441
Lser 2 4 3.819884204E-09
C1 3 4 0.00027
Rpar 3 4 18518.5185185185
.ends 875075355003_270uF
*******
.subckt 875075355004_330uF 1 2
Rser 1 3 0.00891040738169
Lser 2 4 4.040244724E-09
C1 3 4 0.00033
Rpar 3 4 15151.5151515152
.ends 875075355004_330uF
*******
.subckt 875075361005_470uF 1 2
Rser 1 3 0.00824794340995
Lser 2 4 5.241662528E-09
C1 3 4 0.00047
Rpar 3 4 10638.2978723404
.ends 875075361005_470uF
*******
.subckt 875075361006_680uF 1 2
Rser 1 3 0.00907696998223
Lser 2 4 5.257605704E-09
C1 3 4 0.00068
Rpar 3 4 7352.94117647059
.ends 875075361006_680uF
*******
.subckt 875075361007_820uF 1 2
Rser 1 3 0.00783844481106
Lser 2 4 5.11266636E-09
C1 3 4 0.00082
Rpar 3 4 6097.56097560976
.ends 875075361007_820uF
*******
.subckt 875075555001_39uF 1 2
Rser 1 3 0.00894504286591
Lser 2 4 3.860655131E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 875075555001_39uF
*******
.subckt 875075555002_47uF 1 2
Rser 1 3 0.0099786528007
Lser 2 4 4.150163161E-09
C1 3 4 0.000047
Rpar 3 4 106382.978723404
.ends 875075555002_47uF
*******
.subckt 875075555003_68uF 1 2
Rser 1 3 0.0124338939285
Lser 2 4 5.190089124E-09
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 875075555003_68uF
*******
.subckt 875075555004_82uF 1 2
Rser 1 3 0.00958042729986
Lser 2 4 5.09852998E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 875075555004_82uF
*******
.subckt 875075561005_100uF 1 2
Rser 1 3 0.0107963908809
Lser 2 4 7.81186333E-09
C1 3 4 0.0001
Rpar 3 4 50000
.ends 875075561005_100uF
*******
.subckt 875075561006_150uF 1 2
Rser 1 3 0.0118035441314
Lser 2 4 5.709657574E-09
C1 3 4 0.00015
Rpar 3 4 33333.3333333333
.ends 875075561006_150uF
*******
.subckt 875075561007_180uF 1 2
Rser 1 3 0.00884748683423
Lser 2 4 4.968966511E-09
C1 3 4 0.00018
Rpar 3 4 27777.7777777778
.ends 875075561007_180uF
*******
.subckt 875075561008_220uF 1 2
Rser 1 3 0.012154563147
Lser 2 4 5.02464514E-09
C1 3 4 0.00022
Rpar 3 4 22727.2727272727
.ends 875075561008_220uF
*******
.subckt 875075561009_270uF 1 2
Rser 1 3 0.0111482883976
Lser 2 4 5.071280832E-09
C1 3 4 0.00027
Rpar 3 4 18518.5185185185
.ends 875075561009_270uF
*******
.subckt 875075655001_39uF 1 2
Rser 1 3 0.0113149763798
Lser 2 4 5.177745749E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 875075655001_39uF
*******
.subckt 875075655002_68uF 1 2
Rser 1 3 0.01016
Lser 2 4 0.000000003749
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 875075655002_68uF
*******
.subckt 875075655003_82uF 1 2
Rser 1 3 0.00928450836241
Lser 2 4 3.810590877E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 875075655003_82uF
*******
.subckt 875075655005_120uF 1 2
Rser 1 3 0.00974352843849
Lser 2 4 3.790406999E-09
C1 3 4 0.00012
Rpar 3 4 41666.6666666667
.ends 875075655005_120uF
*******
.subckt 875075655006_150uF 1 2
Rser 1 3 0.00946134679851
Lser 2 4 4.074406097E-09
C1 3 4 0.00015
Rpar 3 4 41666.6666666667
.ends 875075655006_150uF
*******
.subckt 875075661004_100uF 1 2
Rser 1 3 0.00860618502417
Lser 2 4 5.47720432E-09
C1 3 4 0.0001
Rpar 3 4 50000
.ends 875075661004_100uF
*******
.subckt 875075661007_180uF 1 2
Rser 1 3 0.0108802573421
Lser 2 4 4.947941742E-09
C1 3 4 0.00018
Rpar 3 4 27777.7777777778
.ends 875075661007_180uF
*******
.subckt 875075661008_220uF 1 2
Rser 1 3 0.0111270909814
Lser 2 4 4.862531768E-09
C1 3 4 0.00022
Rpar 3 4 22727.2727272727
.ends 875075661008_220uF
*******
.subckt 875075661009_270uF 1 2
Rser 1 3 0.0140432856885
Lser 2 4 5.316702808E-09
C1 3 4 0.00027
Rpar 3 4 18518.5185185185
.ends 875075661009_270uF
*******
.subckt 875075661010_330uF 1 2
Rser 1 3 0.0146833185075
Lser 2 4 5.45495338E-09
C1 3 4 0.00033
Rpar 3 4 15151.5151515152
.ends 875075661010_330uF
*******
.subckt 875075755001_10uF 1 2
Rser 1 3 0.0109315812677
Lser 2 4 4.231270383E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 875075755001_10uF
*******
.subckt 875075755002_22uF 1 2
Rser 1 3 0.0140692615854
Lser 2 4 6.022406613E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 875075755002_22uF
*******
.subckt 875075761003_33uF 1 2
Rser 1 3 0.013087585759
Lser 2 4 5.039373348E-09
C1 3 4 0.000033
Rpar 3 4 151515.151515152
.ends 875075761003_33uF
*******
.subckt 875075761004_39uF 1 2
Rser 1 3 0.00858935179083
Lser 2 4 5.45319551E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 875075761004_39uF
*******
.subckt 875075761005_47uF 1 2
Rser 1 3 0.00934111613768
Lser 2 4 5.487187757E-09
C1 3 4 0.000047
Rpar 3 4 106382.978723404
.ends 875075761005_47uF
*******
.subckt 875075761006_56uF 1 2
Rser 1 3 0.0109120399956
Lser 2 4 7.017171452E-09
C1 3 4 0.000056
Rpar 3 4 89285.7142857143
.ends 875075761006_56uF
*******
.subckt 875075761007_68uF 1 2
Rser 1 3 0.0108114773899
Lser 2 4 5.10636587E-09
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 875075761007_68uF
*******
.subckt 875075855001_10uF 1 2
Rser 1 3 0.0108754718643
Lser 2 4 3.969100446E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 875075855001_10uF
*******
.subckt 875075855002_22uF 1 2
Rser 1 3 0.0108615067263
Lser 2 4 4.07194044E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 875075855002_22uF
*******
.subckt 875075855005_39uF 1 2
Rser 1 3 0.0107205858498
Lser 2 4 4.044377124E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 875075855005_39uF
*******
.subckt 875075861003_22uF 1 2
Rser 1 3 0.0091
Lser 2 4 0.000000004
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 875075861003_22uF
*******
.subckt 875075861004_33uF 1 2
Rser 1 3 0.0073
Lser 2 4 0.00000000435
C1 3 4 0.000033
Rpar 3 4 151515.151515152
.ends 875075861004_33uF
*******
.subckt 875075861006_47uF 1 2
Rser 1 3 0.00893031461
Lser 2 4 5.224104755E-09
C1 3 4 0.000047
Rpar 3 4 106382.978723404
.ends 875075861006_47uF
*******
.subckt 875075955001_10uF 1 2
Rser 1 3 0.0143983185003
Lser 2 4 4.173676376E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 875075955001_10uF
*******
.subckt 875075961002_22uF 1 2
Rser 1 3 0.0116062294459
Lser 2 4 5.269169652E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 875075961002_22uF
*******
.subckt 875076155002_12uF 1 2
Rser 1 3 0.0101212388697
Lser 2 4 4.185863478E-09
C1 3 4 0.000012
Rpar 3 4 416666.666666667
.ends 875076155002_12uF
*******
.subckt 875076161003_22uF 1 2
Rser 1 3 0.00882184387393
Lser 2 4 5.398077523E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 875076161003_22uF
*******
