**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ASLI
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         5/31/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 865080140001_22uF 1 2
Rser 1 3 1.4
Lser 2 4 7.03609827E-10
C1 3 4 0.000022
Rpar 3 4 2100000
.ends 865080140001_22uF
*******
.subckt 865080140002_27uF 1 2
Rser 1 3 1.4
Lser 2 4 7.898467596E-09
C1 3 4 0.000027
Rpar 3 4 2100000
.ends 865080140002_27uF
*******
.subckt 865080140003_33uF 1 2
Rser 1 3 1.48
Lser 2 4 0.0000000009785
C1 3 4 0.000033
Rpar 3 4 2100000
.ends 865080140003_33uF
*******
.subckt 865080140004_47uF 1 2
Rser 1 3 1.25
Lser 2 4 0.000000001066
C1 3 4 0.000047
Rpar 3 4 2100000
.ends 865080140004_47uF
*******
.subckt 865080142005_56uF 1 2
Rser 1 3 0.82
Lser 2 4 1.742530489E-09
C1 3 4 0.000056
Rpar 3 4 1784702.54957507
.ends 865080142005_56uF
*******
.subckt 865080142006_68uF 1 2
Rser 1 3 0.704
Lser 2 4 2.37966274140194E-08
C1 3 4 0.000068
Rpar 3 4 1471962.61682243
.ends 865080142006_68uF
*******
.subckt 865080142007_100uF 1 2
Rser 1 3 0.56
Lser 2 4 0.000000002121
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080142007_100uF
*******
.subckt 865080143008_150uF 1 2
Rser 1 3 0.45
Lser 2 4 0.000000002589
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865080143008_150uF
*******
.subckt 865080143009_220uF 1 2
Rser 1 3 0.317
Lser 2 4 2.01727680531737E-08
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080143009_220uF
*******
.subckt 865080145010_330uF 1 2
Rser 1 3 0.177
Lser 2 4 5.56044228297646E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865080145010_330uF
*******
.subckt 865080149011_330uF 1 2
Rser 1 3 0.27
Lser 2 4 0.00000000025
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865080149011_330uF
*******
.subckt 865080153012_470uF 1 2
Rser 1 3 0.132
Lser 2 4 5.14482998700241E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865080153012_470uF
*******
.subckt 865080153013_680uF 1 2
Rser 1 3 0.131
Lser 2 4 6.15086109794052E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865080153013_680uF
*******
.subckt 865080153014_1mF 1 2
Rser 1 3 0.117
Lser 2 4 6.17056298530583E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 865080153014_1mF
*******
.subckt 865080157015_1.2mF 1 2
Rser 1 3 0.134733372703
Lser 2 4 7.519595256E-09
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 865080157015_1.2mF
*******
.subckt 865080157016_1.5mF 1 2
Rser 1 3 0.086
Lser 2 4 7.32576603659146E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 865080157016_1.5mF
*******
.subckt 865080162017_3.3mF 1 2
Rser 1 3 0.0968673260248
Lser 2 4 1.2961682119E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 865080162017_3.3mF
*******
.subckt 865080163018_6.8mF 1 2
Rser 1 3 0.0501343357384
Lser 2 4 1.4162560232E-08
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 865080163018_6.8mF
*******
.subckt 865080240001_22uF 1 2
Rser 1 3 1.4
Lser 2 4 0.00000000105
C1 3 4 0.000022
Rpar 3 4 3333333.33333333
.ends 865080240001_22uF
*******
.subckt 865080240003_33uF 1 2
Rser 1 3 1.36
Lser 2 4 0.000000000864728
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865080240003_33uF
*******
.subckt 865080242002_27uF 1 2
Rser 1 3 1.03
Lser 2 4 0.000000001915
C1 3 4 0.000027
Rpar 3 4 3333333.33333333
.ends 865080242002_27uF
*******
.subckt 865080242004_47uF 1 2
Rser 1 3 0.78
Lser 2 4 0.000000000025
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865080242004_47uF
*******
.subckt 865080243005_56uF 1 2
Rser 1 3 0.56
Lser 2 4 0.000000002444
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 865080243005_56uF
*******
.subckt 865080243006_68uF 1 2
Rser 1 3 0.54
Lser 2 4 0.000000002441
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 865080243006_68uF
*******
.subckt 865080243007_100uF 1 2
Rser 1 3 0.653363834984
Lser 2 4 9.866278783E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080243007_100uF
*******
.subckt 865080243008_150uF 1 2
Rser 1 3 0.45
Lser 2 4 0.000000002592
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865080243008_150uF
*******
.subckt 865080245009_220uF 1 2
Rser 1 3 0.244
Lser 2 4 4.56031232986069E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080245009_220uF
*******
.subckt 865080249010_220uF 1 2
Rser 1 3 0.44328
Lser 2 4 4.089642131E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080249010_220uF
*******
.subckt 865080253011_330uF 1 2
Rser 1 3 0.2305
Lser 2 4 3.888824971E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865080253011_330uF
*******
.subckt 865080253012_470uF 1 2
Rser 1 3 0.14
Lser 2 4 0.0000000006
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865080253012_470uF
*******
.subckt 865080257013_680uF 1 2
Rser 1 3 0.12926
Lser 2 4 5.227999329E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865080257013_680uF
*******
.subckt 865080257014_1mF 1 2
Rser 1 3 0.149063145805
Lser 2 4 7.231052693E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 865080257014_1mF
*******
.subckt 865080262015_2.2mF 1 2
Rser 1 3 0.0919460151431
Lser 2 4 1.1726708153E-08
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 865080262015_2.2mF
*******
.subckt 865080263016_4.7mF 1 2
Rser 1 3 0.046560766426
Lser 2 4 1.7039410182E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 865080263016_4.7mF
*******
.subckt 865080340001_10uF 1 2
Rser 1 3 1.3
Lser 2 4 6.62786597E-10
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 865080340001_10uF
*******
.subckt 865080340002_15uF 1 2
Rser 1 3 1.42
Lser 2 4 0.0000000000023
C1 3 4 0.000015
Rpar 3 4 5333333.33333333
.ends 865080340002_15uF
*******
.subckt 865080340003_22uF 1 2
Rser 1 3 1.48
Lser 2 4 0.000000000971804
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865080340003_22uF
*******
.subckt 865080342004_27uF 1 2
Rser 1 3 0.85
Lser 2 4 0.000000002283
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 865080342004_27uF
*******
.subckt 865080342006_47uF 1 2
Rser 1 3 0.59
Lser 2 4 0.000000000055
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865080342006_47uF
*******
.subckt 865080343005_33uF 1 2
Rser 1 3 0.4
Lser 2 4 0.00000000015
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865080343005_33uF
*******
.subckt 865080343007_56uF 1 2
Rser 1 3 0.6
Lser 2 4 0.000000002347
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 865080343007_56uF
*******
.subckt 865080343008_68uF 1 2
Rser 1 3 0.55
Lser 2 4 0.000000002448
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 865080343008_68uF
*******
.subckt 865080343009_100uF 1 2
Rser 1 3 0.9
Lser 2 4 2.918567665E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080343009_100uF
*******
.subckt 865080345010_150uF 1 2
Rser 1 3 0.42
Lser 2 4 0.000000002527
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865080345010_150uF
*******
.subckt 865080345012_220uF 1 2
Rser 1 3 0.25
Lser 2 4 0.000000002805
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080345012_220uF
*******
.subckt 865080349011_150uF 1 2
Rser 1 3 0.317
Lser 2 4 0.00000000025
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865080349011_150uF
*******
.subckt 865080349013_220uF 1 2
Rser 1 3 0.42719
Lser 2 4 4.405034758E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080349013_220uF
*******
.subckt 865080353014_330uF 1 2
Rser 1 3 0.145
Lser 2 4 0.000000001
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865080353014_330uF
*******
.subckt 865080353015_470uF 1 2
Rser 1 3 0.133
Lser 2 4 2.09657010043051E-08
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865080353015_470uF
*******
.subckt 865080357016_680uF 1 2
Rser 1 3 0.08
Lser 2 4 7.11803919602637E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865080357016_680uF
*******
.subckt 865080362017_1.5mF 1 2
Rser 1 3 0.056
Lser 2 4 8.91133575170173E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 865080362017_1.5mF
*******
.subckt 865080363018_3.3mF 1 2
Rser 1 3 0.0512003095746
Lser 2 4 1.7019727769E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 865080363018_3.3mF
*******
.subckt 865080440001_6.8uF 1 2
Rser 1 3 1.45
Lser 2 4 0.000000000874985
C1 3 4 0.0000068
Rpar 3 4 8333333.33333333
.ends 865080440001_6.8uF
*******
.subckt 865080440002_10uF 1 2
Rser 1 3 1.3
Lser 2 4 6.97769198E-10
C1 3 4 0.00001
Rpar 3 4 8333333.33333333
.ends 865080440002_10uF
*******
.subckt 865080442003_15uF 1 2
Rser 1 3 1.11
Lser 2 4 0.000000001358
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends 865080442003_15uF
*******
.subckt 865080442004_22uF 1 2
Rser 1 3 0.966876169486
Lser 2 4 8.802109939E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865080442004_22uF
*******
.subckt 865080442006_33uF 1 2
Rser 1 3 0.89
Lser 2 4 1.827910305E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865080442006_33uF
*******
.subckt 865080443005_27uF 1 2
Rser 1 3 0.56
Lser 2 4 0.000000002678
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 865080443005_27uF
*******
.subckt 865080443007_47uF 1 2
Rser 1 3 0.39
Lser 2 4 0.000000002583
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865080443007_47uF
*******
.subckt 865080443008_56uF 1 2
Rser 1 3 0.57
Lser 2 4 0.00000000245
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 865080443008_56uF
*******
.subckt 865080443009_68uF 1 2
Rser 1 3 0.43
Lser 2 4 0.000000002866
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 865080443009_68uF
*******
.subckt 865080445010_100uF 1 2
Rser 1 3 0.183
Lser 2 4 4.92952910408854E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080445010_100uF
*******
.subckt 865080449011_100uF 1 2
Rser 1 3 0.284
Lser 2 4 2.1231734564992E-08
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080449011_100uF
*******
.subckt 865080453012_150uF 1 2
Rser 1 3 0.16
Lser 2 4 0.00000000095
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865080453012_150uF
*******
.subckt 865080453013_220uF 1 2
Rser 1 3 0.127
Lser 2 4 5.40044438570286E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080453013_220uF
*******
.subckt 865080453014_330uF 1 2
Rser 1 3 0.1
Lser 2 4 5.94822679517771E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865080453014_330uF
*******
.subckt 865080457015_470uF 1 2
Rser 1 3 0.08
Lser 2 4 0.0000000011
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865080457015_470uF
*******
.subckt 865080462016_1mF 1 2
Rser 1 3 0.0817097292197
Lser 2 4 1.1641816996E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 865080462016_1mF
*******
.subckt 865080463017_2.2mF 1 2
Rser 1 3 0.0509726897787
Lser 2 4 1.3874413766E-08
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 865080463017_2.2mF
*******
.subckt 865080540001_3.3uF 1 2
Rser 1 3 1.03
Lser 2 4 0.000000000016
C1 3 4 0.0000033
Rpar 3 4 11666666.6666667
.ends 865080540001_3.3uF
*******
.subckt 865080540002_4.7uF 1 2
Rser 1 3 1.93954804011
Lser 2 4 1.227468927E-09
C1 3 4 0.0000047
Rpar 3 4 11666666.6666667
.ends 865080540002_4.7uF
*******
.subckt 865080540003_6.8uF 1 2
Rser 1 3 1.4
Lser 2 4 6.37421672E-10
C1 3 4 0.0000068
Rpar 3 4 11666666.6666667
.ends 865080540003_6.8uF
*******
.subckt 865080540004_10uF 1 2
Rser 1 3 1.12
Lser 2 4 0.000000001048
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865080540004_10uF
*******
.subckt 865080542005_15uF 1 2
Rser 1 3 0.89
Lser 2 4 1.787806959E-09
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends 865080542005_15uF
*******
.subckt 865080542006_22uF 1 2
Rser 1 3 0.75
Lser 2 4 0.000000002144
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 865080542006_22uF
*******
.subckt 865080543007_27uF 1 2
Rser 1 3 0.54
Lser 2 4 0.000000002383
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 865080543007_27uF
*******
.subckt 865080543008_33uF 1 2
Rser 1 3 0.355
Lser 2 4 0.00000000022
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865080543008_33uF
*******
.subckt 865080543009_47uF 1 2
Rser 1 3 0.341
Lser 2 4 1.91825309054084E-08
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865080543009_47uF
*******
.subckt 865080545010_56uF 1 2
Rser 1 3 0.34
Lser 2 4 0.000000002667
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 865080545010_56uF
*******
.subckt 865080545011_68uF 1 2
Rser 1 3 0.375
Lser 2 4 0.000000002608
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 865080545011_68uF
*******
.subckt 865080545012_100uF 1 2
Rser 1 3 0.31
Lser 2 4 0.000000002805
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080545012_100uF
*******
.subckt 865080553013_150uF 1 2
Rser 1 3 0.175
Lser 2 4 0.000000001
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865080553013_150uF
*******
.subckt 865080553014_220uF 1 2
Rser 1 3 0.123
Lser 2 4 2.08433561671112E-08
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080553014_220uF
*******
.subckt 865080557015_330uF 1 2
Rser 1 3 0.083
Lser 2 4 0.0000000018
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865080557015_330uF
*******
.subckt 865080562016_470uF 1 2
Rser 1 3 0.0977460160899
Lser 2 4 1.1223380033E-08
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865080562016_470uF
*******
.subckt 865080562017_680uF 1 2
Rser 1 3 0.0782678595762
Lser 2 4 1.0567424615E-08
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 865080562017_680uF
*******
.subckt 865080563018_1.5mF 1 2
Rser 1 3 0.0483494450204
Lser 2 4 1.394324891E-08
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 865080563018_1.5mF
*******
.subckt 865080640001_1uF 1 2
Rser 1 3 2.53014275436
Lser 2 4 1.662056393E-09
C1 3 4 0.000001
Rpar 3 4 16666666.6666667
.ends 865080640001_1uF
*******
.subckt 865080640002_2.2uF 1 2
Rser 1 3 1.67
Lser 2 4 0.000000000594774
C1 3 4 0.0000022
Rpar 3 4 16666666.6666667
.ends 865080640002_2.2uF
*******
.subckt 865080640003_3.3uF 1 2
Rser 1 3 1.86102954548
Lser 2 4 9.72669922E-10
C1 3 4 0.0000033
Rpar 3 4 16666666.6666667
.ends 865080640003_3.3uF
*******
.subckt 865080640004_4.7uF 1 2
Rser 1 3 2.06982211189
Lser 2 4 7.26920671E-10
C1 3 4 0.0000047
Rpar 3 4 16666666.6666667
.ends 865080640004_4.7uF
*******
.subckt 865080642005_6.8uF 1 2
Rser 1 3 1.2
Lser 2 4 0.000000000011
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 865080642005_6.8uF
*******
.subckt 865080642006_10uF 1 2
Rser 1 3 1.18
Lser 2 4 0.000000001208
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865080642006_10uF
*******
.subckt 865080643007_15uF 1 2
Rser 1 3 0.79
Lser 2 4 0.000000002268
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends 865080643007_15uF
*******
.subckt 865080643008_22uF 1 2
Rser 1 3 1.05
Lser 2 4 0.000000002206
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865080643008_22uF
*******
.subckt 865080645009_27uF 1 2
Rser 1 3 0.48
Lser 2 4 0.000000002508
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 865080645009_27uF
*******
.subckt 865080645010_33uF 1 2
Rser 1 3 0.49
Lser 2 4 0.000000002502
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865080645010_33uF
*******
.subckt 865080645012_47uF 1 2
Rser 1 3 0.49
Lser 2 4 0.000000002503
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865080645012_47uF
*******
.subckt 865080649011_33uF 1 2
Rser 1 3 0.64
Lser 2 4 0.000000003917
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865080649011_33uF
*******
.subckt 865080649013_47uF 1 2
Rser 1 3 0.52
Lser 2 4 0.000000003785
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865080649013_47uF
*******
.subckt 865080653014_56uF 1 2
Rser 1 3 0.31
Lser 2 4 0.000000004016
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 865080653014_56uF
*******
.subckt 865080653015_68uF 1 2
Rser 1 3 0.247
Lser 2 4 2.02792396606264E-08
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 865080653015_68uF
*******
.subckt 865080653016_100uF 1 2
Rser 1 3 0.197
Lser 2 4 4.80864427233527E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080653016_100uF
*******
.subckt 865080657017_150uF 1 2
Rser 1 3 0.159
Lser 2 4 2.20414099421022E-08
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865080657017_150uF
*******
.subckt 865080657018_220uF 1 2
Rser 1 3 0.154
Lser 2 4 2.1311583677206E-08
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080657018_220uF
*******
.subckt 865080662019_330uF 1 2
Rser 1 3 0.105
Lser 2 4 2.46796591092533E-08
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865080662019_330uF
*******
.subckt 865080663020_1mF 1 2
Rser 1 3 0.0748540658977
Lser 2 4 1.375834307E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 865080663020_1mF
*******
.subckt 865080740002_100nF 1 2
Rser 1 3 3.18631176928
Lser 2 4 1.586363758E-09
C1 3 4 0.0000001
Rpar 3 4 21000000
.ends 865080740002_100nF
*******
.subckt 865080740003_220nF 1 2
Rser 1 3 1.33746685539
Lser 2 4 1.770799678E-09
C1 3 4 0.00000022
Rpar 3 4 21000000
.ends 865080740003_220nF
*******
.subckt 865080740004_330nF 1 2
Rser 1 3 0.84576
Lser 2 4 1.483085699E-09
C1 3 4 0.00000033
Rpar 3 4 21000000
.ends 865080740004_330nF
*******
.subckt 865080740005_470nF 1 2
Rser 1 3 1.02549967334
Lser 2 4 1.576036423E-09
C1 3 4 0.00000047
Rpar 3 4 21000000
.ends 865080740005_470nF
*******
.subckt 865080740006_1uF 1 2
Rser 1 3 1.14836679496
Lser 2 4 1.843217422E-09
C1 3 4 0.000001
Rpar 3 4 21000000
.ends 865080740006_1uF
*******
.subckt 865080740007_2.2uF 1 2
Rser 1 3 2.6220795198
Lser 2 4 1.245516258E-09
C1 3 4 0.0000022
Rpar 3 4 21000000
.ends 865080740007_2.2uF
*******
.subckt 865080742008_3.3uF 1 2
Rser 1 3 2.26536817678
Lser 2 4 1.632556761E-09
C1 3 4 0.0000033
Rpar 3 4 21000000
.ends 865080742008_3.3uF
*******
.subckt 865080742009_4.7uF 1 2
Rser 1 3 2.01859646658
Lser 2 4 1.319528572E-09
C1 3 4 0.0000047
Rpar 3 4 21000000
.ends 865080742009_4.7uF
*******
.subckt 865080743010_10uF 1 2
Rser 1 3 1.41364915984
Lser 2 4 2.069724096E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865080743010_10uF
*******
.subckt 865080745011_22uF 1 2
Rser 1 3 0.91318
Lser 2 4 2.180712302E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865080745011_22uF
*******
.subckt 865080753012_33uF 1 2
Rser 1 3 0.4
Lser 2 4 3.369105384E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865080753012_33uF
*******
.subckt 865080753013_47uF 1 2
Rser 1 3 0.566
Lser 2 4 3.250953097E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865080753013_47uF
*******
.subckt 865080757014_100uF 1 2
Rser 1 3 0.34505
Lser 2 4 6.070502385E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865080757014_100uF
*******
.subckt 865080762015_220uF 1 2
Rser 1 3 0.12
Lser 2 4 0.000000006344
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865080762015_220uF
*******
.subckt 865080763016_470uF 1 2
Rser 1 3 0.11946
Lser 2 4 2.8524845229E-08
C1 3 4 0.00047
Rpar 3 4 212765.957446808
.ends 865080763016_470uF
*******
.subckt 865080840001_1uF 1 2
Rser 1 3 1.17199906098
Lser 2 4 1.876832606E-09
C1 3 4 0.000001
Rpar 3 4 33333333.3333333
.ends 865080840001_1uF
*******
.subckt 865080843002_2.2uF 1 2
Rser 1 3 1.45580312267
Lser 2 4 2.300919093E-09
C1 3 4 0.0000022
Rpar 3 4 33333333.3333333
.ends 865080843002_2.2uF
*******
.subckt 865080845004_4.7uF 1 2
Rser 1 3 1.20635081633
Lser 2 4 2.429626381E-09
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 865080845004_4.7uF
*******
.subckt 865080845005_10uF 1 2
Rser 1 3 1.22436440935
Lser 2 4 2.282424258E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865080845005_10uF
*******
.subckt 865080853006_22uF 1 2
Rser 1 3 0.921
Lser 2 4 2.802364372E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865080853006_22uF
*******
.subckt 865080857007_33uF 1 2
Rser 1 3 0.014
Lser 2 4 3.006650612E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865080857007_33uF
*******
.subckt 865080862008_47uF 1 2
Rser 1 3 0.363
Lser 2 4 5.766036776E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865080862008_47uF
*******
.subckt 865080863009_150uF 1 2
Rser 1 3 0.25624
Lser 2 4 3.8100112604E-08
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865080863009_150uF
*******
.subckt 865080864003_3.3uF 1 2
Rser 1 3 1.29562227638
Lser 2 4 2.029684343E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 865080864003_3.3uF
*******
.subckt 865081740001_1uF 1 2
Rser 1 3 0.928
Lser 2 4 1.602150004E-09
C1 3 4 0.000001
Rpar 3 4 26666666.6666667
.ends 865081740001_1uF
*******
.subckt 865081742002_2.2uF 1 2
Rser 1 3 1.44253320969
Lser 2 4 1.922620298E-09
C1 3 4 0.0000022
Rpar 3 4 26666666.6666667
.ends 865081742002_2.2uF
*******
.subckt 865081743003_3.3uF 1 2
Rser 1 3 1.23372239357
Lser 2 4 2.210566663E-09
C1 3 4 0.0000033
Rpar 3 4 26666666.6666667
.ends 865081743003_3.3uF
*******
.subckt 865081743004_4.7uF 1 2
Rser 1 3 1.41842773889
Lser 2 4 2.08329908E-09
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 865081743004_4.7uF
*******
.subckt 865081745005_10uF 1 2
Rser 1 3 1.21235944747
Lser 2 4 2.108822089E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865081745005_10uF
*******
.subckt 865081745006_22uF 1 2
Rser 1 3 1.1592262187
Lser 2 4 2.135411412E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 865081745006_22uF
*******
.subckt 865081753007_33uF 1 2
Rser 1 3 0.965
Lser 2 4 2.750209091E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865081753007_33uF
*******
.subckt 865081757008_47uF 1 2
Rser 1 3 0.902
Lser 2 4 5.130649603E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865081757008_47uF
*******
.subckt 865081762009_100uF 1 2
Rser 1 3 0.465
Lser 2 4 5.713520271E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865081762009_100uF
*******
.subckt 865081763010_150uF 1 2
Rser 1 3 0.25064
Lser 2 4 3.605125411E-08
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 865081763010_150uF
*******
.subckt 865081763011_220uF 1 2
Rser 1 3 0.22523
Lser 2 4 2.8406226806E-08
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865081763011_220uF
*******
