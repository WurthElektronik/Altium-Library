**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Coupled Inductor
* Matchcode:              WE-TDC HV 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 8018_76889430056_5.6u  1  2  3  4  PARAMS:
+  Cww=8.6p
+  Rp1=8208
+  Cp1=1.977p
+  Lp1=5.656u
+  Rp2=7955
+  Cp2=1.937p
+  Lp2=5.773u
+  RDC1=0.19
+  RDC2=0.19
+  K=0.976509820007678
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_76889430100_10u  1  2  3  4  PARAMS:
+  Cww=12.4p
+  Rp1=13109
+  Cp1=2.029p
+  Lp1=10.107u
+  Rp2=12977
+  Cp2=1.984p
+  Lp2=10.335u
+  RDC1=0.28
+  RDC2=0.28
+  K=0.983869910099907
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_76889430150_15u  1  2  3  4  PARAMS:
+  Cww=15.2p
+  Rp1=15047
+  Cp1=2.095p
+  Lp1=14.376u
+  Rp2=16822
+  Cp2=2.015p
+  Lp2=14.925u
+  RDC1=0.38
+  RDC2=0.38
+  K=0.986576572463249
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_76889430220_22u  1  2  3  4  PARAMS:
+  Cww=17.8p
+  Rp1=21154
+  Cp1=1.94p
+  Lp1=23.731u
+  Rp2=22726
+  Cp2=1.925p
+  Lp2=23.91u
+  RDC1=0.7
+  RDC2=0.7
+  K=0.983962305264698
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_76889440047_4.7u  1  2  3  4  PARAMS:
+  Cww=12.6p
+  Rp1=7500
+  Cp1=3.185p
+  Lp1=4.296u
+  Rp2=6917
+  Cp2=3.174p
+  Lp2=4.312u
+  RDC1=0.085
+  RDC2=0.085
+  K=0.987151500584578
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_76889440100_10u  1  2  3  4  PARAMS:
+  Cww=24.3p
+  Rp1=9559
+  Cp1=3.858p
+  Lp1=9.541u
+  Rp2=8982
+  Cp2=3.914p
+  Lp2=9.583u
+  RDC1=0.16
+  RDC2=0.16
+  K=0.986407623652615
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_76889440150_15u  1  2  3  4  PARAMS:
+  Cww=25.9p
+  Rp1=18540
+  Cp1=3.658p
+  Lp1=15.397u
+  Rp2=17890
+  Cp2=3.697p
+  Lp2=15.234u
+  RDC1=0.3
+  RDC2=0.3
+  K=0.987252078583108
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_76889440220_22u  1  2  3  4  PARAMS:
+  Cww=26.4p
+  Rp1=22949
+  Cp1=4.049p
+  Lp1=20.842u
+  Rp2=25003
+  Cp2=4.096p
+  Lp2=20.599u
+  RDC1=0.39
+  RDC2=0.39
+  K=0.987420882906575
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_76889440330_33u  1  2  3  4  PARAMS:
+  Cww=28.5p
+  Rp1=25849
+  Cp1=4.343p
+  Lp1=35.633u
+  Rp2=25432
+  Cp2=4.343p
+  Lp2=35.63u
+  RDC1=0.575
+  RDC2=0.575
+  K=0.990102535247249
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
