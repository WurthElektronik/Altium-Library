**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Shielded Power Inductor
* Matchcode:             WE-XHMI
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         5/13/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1090_74439369015_1.5u 1 2
Rp 1 2 1195
Cp 1 2 19.206p
Rs 1 N3 0.00146
L1 N3 2 1.349u
.ends 1090_74439369015_1.5u
*******
.subckt 1090_74439369022_2.2u 1 2
Rp 1 2 2074
Cp 1 2 14.601p
Rs 1 N3 0.0022
L1 N3 2 2.242u
.ends 1090_74439369022_2.2u
*******
.subckt 1090_74439369033_3.3u 1 2
Rp 1 2 3017
Cp 1 2 14.697p
Rs 1 N3 0.0034
L1 N3 2 3.164u
.ends 1090_74439369033_3.3u
*******
.subckt 1090_74439369047_4.7u 1 2
Rp 1 2 4114
Cp 1 2 12.704p
Rs 1 N3 0.005
L1 N3 2 4.625u
.ends 1090_74439369047_4.7u
*******
.subckt 1090_74439369056_5.6u 1 2
Rp 1 2 4898
Cp 1 2 13.52p
Rs 1 N3 0.0059
L1 N3 2 5.491u
.ends 1090_74439369056_5.6u
*******
.subckt 1090_74439369068_6.8u 1 2
Rp 1 2 5791
Cp 1 2 14.891p
Rs 1 N3 0.00716
L1 N3 2 7.08u
.ends 1090_74439369068_6.8u
*******
.subckt 1090_74439369082_8.2u 1 2
Rp 1 2 7214
Cp 1 2 12.059p
Rs 1 N3 0.01
L1 N3 2 8.743u
.ends 1090_74439369082_8.2u
*******
.subckt 1090_74439369100_10u 1 2
Rp 1 2 7876
Cp 1 2 13.203p
Rs 1 N3 0.011
L1 N3 2 10.09u
.ends 1090_74439369100_10u
*******
.subckt 1090_74439369150_15u 1 2
Rp 1 2 8204
Cp 1 2 14.622p
Rs 1 N3 0.0148
L1 N3 2 14.546u
.ends 1090_74439369150_15u
*******
.subckt 1510_74439370047_4.7u 1 2
Rp 1 2 4296
Cp 1 2 22.242p
Rs 1 N3 0.0031
L1 N3 2 4.217u
.ends 1510_74439370047_4.7u
*******
.subckt 1510_74439370068_6.8u 1 2
Rp 1 2 5066
Cp 1 2 21.801p
Rs 1 N3 0.0041
L1 N3 2 6.111u
.ends 1510_74439370068_6.8u
*******
.subckt 1510_74439370082_8.2u 1 2
Rp 1 2 6284
Cp 1 2 25.54p
Rs 1 N3 0.0055
L1 N3 2 8.328u
.ends 1510_74439370082_8.2u
*******
.subckt 1510_74439370100_10u 1 2
Rp 1 2 5244
Cp 1 2 29.045p
Rs 1 N3 0.0064
L1 N3 2 10.4u
.ends 1510_74439370100_10u
*******
.subckt 1510_74439370150_15u 1 2
Rp 1 2 7827
Cp 1 2 24.013p
Rs 1 N3 0.0105
L1 N3 2 15.895u
.ends 1510_74439370150_15u
*******
.subckt 1510_74439370220_22u 1 2
Rp 1 2 8204
Cp 1 2 26.195p
Rs 1 N3 0.0125
L1 N3 2 20.695u
.ends 1510_74439370220_22u
*******
.subckt 1510_74439370330_33u 1 2
Rp 1 2 10776
Cp 1 2 27.127p
Rs 1 N3 0.018
L1 N3 2 31.904u
.ends 1510_74439370330_33u
*******
.subckt 6030_744393440015_0.15u 1 2
Rp 1 2 306.09
Cp 1 2 4.722p
Rs 1 N3 0.00124
L1 N3 2 0.147u
.ends 6030_744393440015_0.15u
*******
.subckt 6030_744393440018_0.18u 1 2
Rp 1 2 393.041
Cp 1 2 5.062p
Rs 1 N3 0.00132
L1 N3 2 0.176u
.ends 6030_744393440018_0.18u
*******
.subckt 6030_744393440033_0.33u 1 2
Rp 1 2 683.781
Cp 1 2 6.324p
Rs 1 N3 0.0021
L1 N3 2 0.316u
.ends 6030_744393440033_0.33u
*******
.subckt 6030_744393440056_0.56u 1 2
Rp 1 2 876.79
Cp 1 2 7.515p
Rs 1 N3 0.0029
L1 N3 2 0.561u
.ends 6030_744393440056_0.56u
*******
.subckt 6030_74439344010_1u 1 2
Rp 1 2 1956
Cp 1 2 7.102p
Rs 1 N3 0.0055
L1 N3 2 1.008u
.ends 6030_74439344010_1u
*******
.subckt 6030_74439344012_1.2u 1 2
Rp 1 2 2178
Cp 1 2 8.182p
Rs 1 N3 0.0064
L1 N3 2 1.105u
.ends 6030_74439344012_1.2u
*******
.subckt 6030_74439344022_2.2u 1 2
Rp 1 2 2927
Cp 1 2 8.36p
Rs 1 N3 0.0105
L1 N3 2 2.182u
.ends 6030_74439344022_2.2u
*******
.subckt 6030_74439344033_3.3u 1 2
Rp 1 2 4970
Cp 1 2 7.979p
Rs 1 N3 0.0192
L1 N3 2 3.247u
.ends 6030_74439344033_3.3u
*******
.subckt 6030_74439344047_4.7u 1 2
Rp 1 2 7211
Cp 1 2 7.002p
Rs 1 N3 0.031
L1 N3 2 4.676u
.ends 6030_74439344047_4.7u
*******
.subckt 6060_74439346010_1u 1 2
Rp 1 2 1210
Cp 1 2 6.845p
Rs 1 N3 0.00339
L1 N3 2 1.046u
.ends 6060_74439346010_1u
*******
.subckt 6060_74439346012_1.2u 1 2
Rp 1 2 1330
Cp 1 2 8.78p
Rs 1 N3 0.00365
L1 N3 2 1.158u
.ends 6060_74439346012_1.2u
*******
.subckt 6060_74439346015_1.5u 1 2
Rp 1 2 1396
Cp 1 2 9.359p
Rs 1 N3 0.0039
L1 N3 2 1.373u
.ends 6060_74439346015_1.5u
*******
.subckt 6060_74439346018_1.8u 1 2
Rp 1 2 1659
Cp 1 2 7.994p
Rs 1 N3 0.0047
L1 N3 2 1.806u
.ends 6060_74439346018_1.8u
*******
.subckt 6060_74439346022_2.2u 1 2
Rp 1 2 1877
Cp 1 2 8.362p
Rs 1 N3 0.00558
L1 N3 2 2.182u
.ends 6060_74439346022_2.2u
*******
.subckt 6060_74439346033_3.3u 1 2
Rp 1 2 2955
Cp 1 2 8.785p
Rs 1 N3 0.01083
L1 N3 2 2.95u
.ends 6060_74439346033_3.3u
*******
.subckt 6060_74439346047_4.7u 1 2
Rp 1 2 4305
Cp 1 2 7.633p
Rs 1 N3 0.013
L1 N3 2 4.289u
.ends 6060_74439346047_4.7u
*******
.subckt 6060_74439346056_5.6u 1 2
Rp 1 2 5112
Cp 1 2 7.79p
Rs 1 N3 0.015
L1 N3 2 5.311u
.ends 6060_74439346056_5.6u
*******
.subckt 6060_74439346068_6.8u 1 2
Rp 1 2 5867
Cp 1 2 7.976p
Rs 1 N3 0.0176
L1 N3 2 6.553u
.ends 6060_74439346068_6.8u
*******
.subckt 6060_74439346082_8.2u 1 2
Rp 1 2 6820
Cp 1 2 8.668p
Rs 1 N3 0.023
L1 N3 2 7.855u
.ends 6060_74439346082_8.2u
*******
.subckt 6060_74439346100_10u 1 2
Rp 1 2 9786
Cp 1 2 8.192p
Rs 1 N3 0.0265
L1 N3 2 9.539u
.ends 6060_74439346100_10u
*******
.subckt 6060_74439346150_15u 1 2
Rp 1 2 11178
Cp 1 2 8.829p
Rs 1 N3 0.042
L1 N3 2 15.089u
.ends 6060_74439346150_15u
*******
.subckt 8080_744393580068_0.68u 1 2
Rp 1 2 1027
Cp 1 2 9.182p
Rs 1 N3 0.00141
L1 N3 2 0.71u
.ends 8080_744393580068_0.68u
*******
.subckt 8080_74439358010_1u 1 2
Rp 1 2 1445
Cp 1 2 8.916p
Rs 1 N3 0.0021
L1 N3 2 1.014u
.ends 8080_74439358010_1u
*******
.subckt 8080_74439358015_1.5u 1 2
Rp 1 2 1599
Cp 1 2 11.49p
Rs 1 N3 0.00291
L1 N3 2 1.588u
.ends 8080_74439358015_1.5u
*******
.subckt 8080_74439358022_2.2u 1 2
Rp 1 2 2282
Cp 1 2 10.434p
Rs 1 N3 0.0037
L1 N3 2 2.209u
.ends 8080_74439358022_2.2u
*******
.subckt 8080_74439358047_4.7u 1 2
Rp 1 2 4439
Cp 1 2 10.924p
Rs 1 N3 0.00865
L1 N3 2 4.785u
.ends 8080_74439358047_4.7u
*******
.subckt 8080_74439358068_6.8u 1 2
Rp 1 2 6545
Cp 1 2 7.924p
Rs 1 N3 0.013
L1 N3 2 6.596u
.ends 8080_74439358068_6.8u
*******
.subckt 8080_74439358100_10u 1 2
Rp 1 2 8417
Cp 1 2 8.116p
Rs 1 N3 0.019
L1 N3 2 10.282u
.ends 8080_74439358100_10u
*******
.subckt 8080_74439358150_15u 1 2
Rp 1 2 8485
Cp 1 2 11.885p
Rs 1 N3 0.025
L1 N3 2 14.163u
.ends 8080_74439358150_15u
*******
