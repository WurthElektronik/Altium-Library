**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Molded Coupled Inductor 
* Matchcode:              WE-MCRI
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1090_7448990010_1u  1  2  3  4  PARAMS:
+  Cww=76p
+  Rp1=2131
+  Cp1=18.45p
+  Lp1=1.112u
+  Rp2=2113
+  Cp2=19.055p
+  Lp2=1.076u
+  RDC1=0.007
+  RDC2=0.007
+  K=0.9
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990015_1.5u  1  2  3  4  PARAMS:
+  Cww=79p
+  Rp1=2700
+  Cp1=19.49p
+  Lp1=1.454u
+  Rp2=2741
+  Cp2=19.35p
+  Lp2=1.554u
+  RDC1=0.016
+  RDC2=0.016
+  K=0.921592824046137
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990022_2.2u  1  2  3  4  PARAMS:
+  Cww=90p
+  Rp1=4880
+  Cp1=26.707p
+  Lp1=2.555u
+  Rp2=4518
+  Cp2=26.989p
+  Lp2=2.528u
+  RDC1=0.022
+  RDC2=0.022
+  K=0.945082968940727
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990033_3.3u  1  2  3  4  PARAMS:
+  Cww=99p
+  Rp1=6700
+  Cp1=20.581p
+  Lp1=3.316u
+  Rp2=6635
+  Cp2=20.7p
+  Lp2=3.297u
+  RDC1=0.028
+  RDC2=0.028
+  K=0.9613752775282
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990047_4.7u  1  2  3  4  PARAMS:
+  Cww=98p
+  Rp1=4913
+  Cp1=22.582p
+  Lp1=4.574u
+  Rp2=5004
+  Cp2=22.507p
+  Lp2=4.559u
+  RDC1=0.035
+  RDC2=0.035
+  K=0.972275243403929
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990068_6.8u  1  2  3  4  PARAMS:
+  Cww=131p
+  Rp1=6400
+  Cp1=23.196p
+  Lp1=6.671u
+  Rp2=6631
+  Cp2=23.057p
+  Lp2=6.712u
+  RDC1=0.048
+  RDC2=0.048
+  K=0.980696031338127
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990082_8.2u  1  2  3  4  PARAMS:
+  Cww=162p
+  Rp1=4896
+  Cp1=25.504p
+  Lp1=8.998u
+  Rp2=4972
+  Cp2=25.148p
+  Lp2=9.125u
+  RDC1=0.059
+  RDC2=0.059
+  K=0.983398785199426
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990100_10u  1  2  3  4  PARAMS:
+  Cww=178p
+  Rp1=7321
+  Cp1=28.172p
+  Lp1=10.072u
+  Rp2=7421
+  Cp2=28.127p
+  Lp2=10.088u
+  RDC1=0.064
+  RDC2=0.064
+  K=0.986154146165801
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990150_15u  1  2  3  4  PARAMS:
+  Cww=199p
+  Rp1=8298
+  Cp1=26.456p
+  Lp1=15.755u
+  Rp2=8175
+  Cp2=26.386p
+  Lp2=15.757u
+  RDC1=0.075
+  RDC2=0.075
+  K=0.990252493054171
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990220_22u  1  2  3  4  PARAMS:
+  Cww=226p
+  Rp1=9865
+  Cp1=24.449p
+  Lp1=20.839u
+  Rp2=10350
+  Cp2=24.482p
+  Lp2=20.811u
+  RDC1=0.099
+  RDC2=0.099
+  K=0.99304398877208
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990330_33u  1  2  3  4  PARAMS:
+  Cww=345p
+  Rp1=11110
+  Cp1=29.2p
+  Lp1=32.34u
+  Rp2=11322
+  Cp2=29.225p
+  Lp2=32.429u
+  RDC1=0.129
+  RDC2=0.129
+  K=0.994530496812898
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 1090_7448990470_47u  1  2  3  4  PARAMS:
+  Cww=363p
+  Rp1=26460
+  Cp1=26.452p
+  Lp1=44.153u
+  Rp2=28240
+  Cp2=29.49p
+  Lp2=44.089u
+  RDC1=0.222
+  RDC2=0.222
+  K=0.996162850909386
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
