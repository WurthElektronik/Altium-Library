**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Full-color Top LED Diffused 
* Matchcode:              WL-SFTD
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-17
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1616_150161M153130 1 2 3 4 
D1 1 2 Red
.MODEL Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
D2 1 3 Green
.MODEL Green D
+ IS=75.763E-18
+ N=3.3919
+ RS=.54629
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
D3 1 4 Blue
.MODEL Blue D
+ IS=150.13E-18
+ N=3.3919
+ RS=.5463
+ IKF=413.18E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
.ends
*****************
.subckt 2022_150202M153130 1 2 3 4 
D1 1 2 Red
.MODEL Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
D2 1 3 Green
.MODEL Green D
+ IS=75.763E-18
+ N=3.3919
+ RS=.54629
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
D3 1 4 Blue
.MODEL Blue D
+ IS=150.13E-18
+ N=3.3919
+ RS=.5463
+ IKF=413.18E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
.ends
*****************
.subckt 2828_150282M153310 1 2 3 4 5 6
D1 4 3 Blue
.MODEL Blue D
+ IS=150.13E-18
+ N=3.3919
+ RS=.5463
+ IKF=413.18E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
D2 5 2 Green
.MODEL Green D
+ IS=75.763E-18
+ N=3.3919
+ RS=.54629
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
D3 6 1 Red
.MODEL Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
.ends
*****************
.subckt 3535_150353M153300 1 2 3 4 5 6
D1 1 2 Red
.MODEL Red D
+ IS=843.65E-18
+ N=2.3334
+ RS=.35062
+ IKF=755.09E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
D2 3 4 Green
.MODEL Green D
+ IS=17.287E-12
+ N=4.9970
+ RS=1.9544
+ IKF=356.06E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
D3 5 6 Blue
.MODEL Blue D
+ IS=488.35E-12
+ N=4.4633
+ RS=1.5487
+ IKF=779.60E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=6.00E-6
+ TT=5.0000E-9
.ends
*****************

































