**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Thinfilm Chip Inductor 
* Matchcode:              WE-TCI 
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Ella      
* Date and Time:          2022-06-22
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0201_744900010_1n 1 2
C1 1 N7 320.3197f
L1 1 N1 0.95n
L2 N1 N2 84.0495p
L3 N2 N3 34.6674p
L4 N3 N4 280.2628p
L5 N4 N5 78.4955p
L6 N5 N6 56.0008p
R1 2 N1 868.7166m
R2 2 N2 747.7590m
R3 2 N3 297.4903m
R4 2 N4 561.8773m
R5 2 N5 562.7613m
R6 2 N6 225.3587m
R7 2 N7 2.5725
R8 2 1 10g
.ends 
*******
.subckt 0201_744900012_1.2n 1 2
C1 1 N7 142.2417f
L1 1 N1 1.15n
L2 N1 N2 90.8090p
L3 N2 N3 64.7608p
L4 N3 N4 335.8757p
L5 N4 N5 78.7053p
L6 N5 N6 56.0762p
R1 2 N1 828.9126m
R2 2 N2 769.8246m
R3 2 N3 399.8134m
R4 2 N4 561.0837m
R5 2 N5 558.7898m
R6 2 N6 225.0624m
R7 2 N7 2.5718
R8 2 1 10g
.ends 
*******
.subckt 0201_744900013_1.3n 1 2
C1 1 N7 140.5520f
L1 1 N1 1.25n
L2 N1 N2 93.1279p
L3 N2 N3 40.1304p
L4 N3 N4 280.3138p
L5 N4 N5 78.4954p
L6 N5 N6 56.0008p
R1 2 N1 869.0054m
R2 2 N2 748.0864m
R3 2 N3 298.4877m
R4 2 N4 561.8953m
R5 2 N5 562.7780m
R6 2 N6 225.3598m
R7 2 N7 2.5725
R8 2 1 10g
.ends 
*******
.subckt 0201_744900014_1.4n 1 2
C1 1 N7 223.37f
L1 1 N1 1.33n
L2 N1 N2 98.4726p
L3 N2 N3 46.4725p
L4 N3 N4 280.7142p
L5 N4 N5 78.4970p
L6 N5 N6 56.0017p
R1 2 N1 868.6413m
R2 2 N2 748.5286m
R3 2 N3 300.7126m
R4 2 N4 562.0245m
R5 2 N5 562.8900m
R6 2 N6 225.3664m
R7 2 N7 2.5725
R8 2 1 10g
.ends 
*******
.subckt 0201_744900015_1.5n 1 2
C1 1 N7 208.48f
L1 1 N1 1.43n
L2 N1 N2 110.3201p
L3 N2 N3 55.6799p
L4 N3 N4 344.0937p
L5 N4 N5 78.8777p
L6 N5 N6 56.2099p
R1 2 N1 951.9239m
R2 2 N2 770.0270m
R3 2 N3 419.4204m
R4 2 N4 583.5672m
R5 2 N5 581.6298m
R6 2 N6 226.4618m
R7 2 N7 2.5769
R8 2 1 10g
.ends 
*******
.subckt 0201_744900018_1.8n 1 2
C1 1 N7 173.73f
L1 1 N1 1.7n
L2 N1 N2 143.9246p
L3 N2 N3 216.0225p
L4 N3 N4 208.5669p
L5 N4 N5 8.3803p
L6 N5 N6 37.7011p
R1 2 N1 5.633
R2 2 N2 610.2852m
R3 2 N3 3.559
R4 2 N4 3.9329
R5 2 N5 3.1801
R6 2 N6 3.2396
R7 2 N7 2.6351
R8 2 1 10g
.ends 
*******
.subckt 0201_744900019_1.9n 1 2
C1 1 N7 164.589f
L1 1 N1 1.82n
L2 N1 N2 163.5430p
L3 N2 N3 257.2243p
L4 N3 N4 225.1563p
L5 N4 N5 8.4486p
L6 N5 N6 37.7234p
R1 2 N1 5.6322
R2 2 N2 695.6538m
R3 2 N3 3.5599
R4 2 N4 3.9328
R5 2 N5 3.18
R6 2 N6 3.2395
R7 2 N7 2.6351
R8 2 1 10g
.ends 
*******
.subckt 0201_744900020_2n 1 2
C1 1 N7 200f
L1 1 N1 1.9n
L2 N1 N2 220.1397p
L3 N2 N3 502.4286p
L4 N3 N4 323.8605p
L5 N4 N5 8.9573p
L6 N5 N6 37.8416p
R1 2 N1 5.6212
R2 2 N2 1.1154
R3 2 N3 3.5649
R4 2 N4 3.9311
R5 2 N5 3.1772
R6 2 N6 3.2365
R7 2 N7 2.6351
R8 2 1 10g
.ends 
*******
.subckt 0201_744900022_2.2n 1 2
C1 1 N7 179.5657f
L1 1 N1 2.1n
L2 N1 N2 195.7870p
L3 N2 N3 319.9084p
L4 N3 N4 240.1134p
L5 N4 N5 8.5208p
L6 N5 N6 37.7367p
R1 2 N1 3.1137
R2 2 N2 812.1823m
R3 2 N3 3.253
R4 2 N4 2.9269
R5 2 N5 3.1711
R6 2 N6 3.2309
R7 2 N7 2.5351
R8 2 1 10g
.ends 
*******
.subckt 0201_744900027_2.7n 1 2
C1 1 N7 148.9275f
L1 1 N1 2.5n
L2 N1 N2 322.5951p
L3 N2 N3 796.0514p
L4 N3 N4 484.3178p
L5 N4 N5 9.5766p
L6 N5 N6 37.9918p
R1 2 N1 3.0218
R2 2 N2 1.491
R3 2 N3 3.2863
R4 2 N4 2.9461
R5 2 N5 3.1871
R6 2 N6 3.2457
R7 2 N7 2.535
R8 2 1 10g
.ends 
*******
.subckt 0201_744900033_3.3n 1 2
C1 1 N7 219.4097f
L1 1 N1 3.1n
L2 N1 N2 241.6207p
L3 N2 N3 125.2954p
L4 N3 N4 421.3842p
L5 N4 N5 78.9649p
L6 N5 N6 56.3831p
R1 2 N1 1.9487
R2 2 N2 1.6071
R3 2 N3 1.1745
R4 2 N4 567.7369m
R5 2 N5 564.5155m
R6 2 N6 254.0190m
R7 2 N7 2.5433
R8 2 1 10g
.ends 
*******
.subckt 0201_744900039_3.9n 1 2
C1 1 N7 200.1322f
L1 1 N1 3.65n
L2 N1 N2 380.9044p
L3 N2 N3 186.0649p
L4 N3 N4 2.0982n
L5 N4 N5 87.3919p
L6 N5 N6 59.1879p
R1 2 N1 2.6995
R2 2 N2 2.3471
R3 2 N3 1.6353
R4 2 N4 1.679
R5 2 N5 1.6776
R6 2 N6 1.6636
R7 2 N7 2.5206
R8 2 1 10g
.ends 
*******
.subckt 0201_744900047_4.7n 1 2
C1 1 N7 178.4124f
L1 1 N1 4.4n
L2 N1 N2 458.2869p
L3 N2 N3 224.4762p
L4 N3 N4 1.0824n
L5 N4 N5 82.5216p
L6 N5 N6 57.7641p
R1 2 N1 2.8434
R2 2 N2 2.4959
R3 2 N3 1.3067
R4 2 N4 1.3487
R5 2 N5 1.3754
R6 2 N6 1.3655
R7 2 N7 2.5098
R8 2 1 10g
.ends 
*******
.subckt 0201_744900056_5.6n 1 2
C1 1 N7 241.0831f
L1 1 N1 5.2n
L2 N1 N2 46.4887p
L3 N2 N3 730.2516p
L4 N3 N4 1.5904n
L5 N4 N5 104.9129p
L6 N5 N6 64.7120p
R1 2 N1 11.5022
R2 2 N2 5.2127
R3 2 N3 6.2217
R4 2 N4 4.5263
R5 2 N5 4.4849
R6 2 N6 4.4667
R7 2 N7 4.6411
R8 2 1 10g
.ends 
*******
.subckt 0201_744900068_6.8n 1 2
C1 1 N7 239.5178f
L1 1 N1 6.42n
L2 N1 N2 841.1355p
L3 N2 N3 892.7727p
L4 N3 N4 17.6672n
L5 N4 N5 86.3824p
L6 N5 N6 59.0931p
R1 2 N1 2.8797
R2 2 N2 2.5438
R3 2 N3 982.1425m
R4 2 N4 3.6552
R5 2 N5 3.6779
R6 2 N6 3.7180
R7 2 N7 2.7618
R8 2 1 10g
.ends 
*******
.subckt 0201_744900082_8.2n 1 2
C1 1 N7 221.0935f
L1 1 N1 7.6n
L2 N1 N2 1.3608n
L3 N2 N3 535.6902p
L4 N3 N4 18.3393n
L5 N4 N5 87.9997p
L6 N5 N6 60.8787p
R1 2 N1 4.0745
R2 2 N2 2.6895
R3 2 N3 1.6358
R4 2 N4 2.8266
R5 2 N5 2.8214
R6 2 N6 2.8170
R7 2 N7 2.7866
R8 2 1 10g
.ends 
*******
.subckt 0201_744900110_10n 1 2
C1 1 N7 205.5229f
L1 1 N1 9.3n
L2 N1 N2 1.2335n
L3 N2 N3 1.0514n
L4 N3 N4 110.5220p
L5 N4 N5 96.4875p
L6 N5 N6 62.0536p
R1 2 N1 5.8268
R2 2 N2 3.2525
R3 2 N3 4.8885
R4 2 N4 2.8068
R5 2 N5 2.7748
R6 2 N6 2.7592
R7 2 N7 5.4977
R8 2 1 10g
.ends 
*******
.subckt 0402_744901010_1n 1 2
C1 1 N7 137.4402f
L1 1 N1 0.97n
L2 N1 N2 52.4201p
L3 N2 N3 27.2408p
L4 N3 N4 103.7710p
L5 N4 N5 77.2573p
L6 N5 N6 55.3388p
R1 2 N1 483.4069m
R2 2 N2 373.1065m
R3 2 N3 222.6287m
R4 2 N4 238.4874m
R5 2 N5 149.4495m
R6 2 N6 145.7099m
R7 2 N7 2.1699
R8 2 1 10g
.ends 
*******
.subckt 0402_744901012_1.2n 1 2
C1 1 N7 138.5104f
L1 1 N1 1.15n
L2 N1 N2 89.2053p
L3 N2 N3 45.8128p
L4 N3 N4 458.4447p
L5 N4 N5 78.9395p
L6 N5 N6 55.8111p
R1 2 N1 789.9339m
R2 2 N2 628.2599m
R3 2 N3 531.2235m
R4 2 N4 459.7557m
R5 2 N5 314.2502m
R6 2 N6 302.2874m
R7 2 N7 2.3695
R8 2 1 10g
.ends 
*******
.subckt 0402_744901015_1.5n 1 2
C1 1 N7 168.6589f
L1 1 N1 1.45n
L2 N1 N2 88.8579p
L3 N2 N3 43.7178p
L4 N3 N4 359.6747p
L5 N4 N5 78.5189p
L6 N5 N6 55.7212p
R1 2 N1 726.2627m
R2 2 N2 556.5536m
R3 2 N3 427.7572m
R4 2 N4 349.2647m
R5 2 N5 306.7484m
R6 2 N6 297.7737m
R7 2 N7 2.17
R8 2 1 10g
.ends 
*******
.subckt 0402_744901018_1.8n 1 2
C1 1 N7 241.3279f
L1 1 N1 1.72n
L2 N1 N2 95.5050p
L3 N2 N3 45.2070p
L4 N3 N4 357.0530p
L5 N4 N5 78.5154p
L6 N5 N6 55.7313p
R1 2 N1 803.4264m
R2 2 N2 584.9767m
R3 2 N3 436.9148m
R4 2 N4 349.3554m
R5 2 N5 307.2919m
R6 2 N6 298.4366m
R7 2 N7 2.1707
R8 2 1 10g
.ends 
*******
.subckt 0402_744901022_2.2n 1 2
C1 1 N7 105.1046f
L1 1 N1 2.1n
L2 N1 N2 99.0509p
L3 N2 N3 71.1298p
L4 N3 N4 294.3856p
L5 N4 N5 79.6615p
L6 N5 N6 56.3710p
R1 2 N1 1.7784
R2 2 N2 772.0033m
R3 2 N3 655.6709m
R4 2 N4 377.3181m
R5 2 N5 346.7527m
R6 2 N6 335.3020m
R7 2 N7 2.1639
R8 2 1 10g
.ends 
*******
.subckt 0402_744901027_2.7n 1 2
C1 1 N7 158.2310f
L1 1 N1 2.6n
L2 N1 N2 118.2381p
L3 N2 N3 77.6251p
L4 N3 N4 362.1417p
L5 N4 N5 79.9865p
L6 N5 N6 56.4821p
R1 2 N1 1.7989
R2 2 N2 900.1240m
R3 2 N3 713.4635m
R4 2 N4 398.7051m
R5 2 N5 365.9345m
R6 2 N6 353.0908m
R7 2 N7 2.1641
R8 2 1 10g
.ends 
*******
.subckt 0402_744901030_3n 1 2
C1 1 N7 245.0860f
L1 1 N1 2.85n
L2 N1 N2 135.0696p
L3 N2 N3 83.1800p
L4 N3 N4 302.4298p
L5 N4 N5 79.7336p
L6 N5 N6 56.4619p
R1 2 N1 970.2580m
R2 2 N2 644.7486m
R3 2 N3 564.9297m
R4 2 N4 299.9820m
R5 2 N5 252.6577m
R6 2 N6 228.9269m
R7 2 N7 1.8623
R8 2 1 10g
.ends 
*******
.subckt 0402_744901033_3.3n 1 2
C1 1 N7 219.6216f
L1 1 N1 3.1n
L2 N1 N2 182.8161p
L3 N2 N3 99.6211p
L4 N3 N4 553.9172p
L5 N4 N5 80.9225p
L6 N5 N6 56.8204p
R1 2 N1 1.3498
R2 2 N2 1.0302
R3 2 N3 775.9617m
R4 2 N4 412.9306m
R5 2 N5 372.5798m
R6 2 N6 355.0566m
R7 2 N7 1.8457
R8 2 1 10g
.ends 
*******
.subckt 0402_744901036_3.6n 1 2
C1 1 N7 294.2650f
L1 1 N1 3.4n
L2 N1 N2 297.8214p
L3 N2 N3 340.6494p
L4 N3 N4 407.0730p
L5 N4 N5 343.6793p
L6 N5 N6 72.0079p
R1 2 N1 1.2397
R2 2 N2 358.5687m
R3 2 N3 165.6011m
R4 2 N4 203.2069m
R5 2 N5 130.2723m
R6 2 N6 47.8864m
R7 2 N7 1.9181
R8 2 1 10g
.ends 
*******
.subckt 0402_744901039_3.9n 1 2
C1 1 N7 210.3776f
L1 1 N1 3.6n
L2 N1 N2 310.5648p
L3 N2 N3 100.6399p
L4 N3 N4 634.8364p
L5 N4 N5 78.9111p
L6 N5 N6 56.5082p
R1 2 N1 1.3557
R2 2 N2 1.0496
R3 2 N3 805.8332m
R4 2 N4 459.8370m
R5 2 N5 421.7908m
R6 2 N6 405.6598m
R7 2 N7 1.8461
R8 2 1 10g
.ends 
*******
.subckt 0402_744901043_4.3n 1 2
C1 1 N7 160f
L1 1 N1 4n
L2 N1 N2 337.8586p
L3 N2 N3 103.2687p
L4 N3 N4 964.7055p
L5 N4 N5 80.5879p
L6 N5 N6 57.0135p
R1 2 N1 1.1107
R2 2 N2 822.2528m
R3 2 N3 945.0814m
R4 2 N4 666.3023m
R5 2 N5 635.3236m
R6 2 N6 623.1158m
R7 2 N7 1.6469
R8 2 1 10g
.ends 
*******
.subckt 0402_744901047_4.7n 1 2
C1 1 N7 138.4383f
L1 1 N1 4.4n
L2 N1 N2 270.4757p
L3 N2 N3 103.2200p
L4 N3 N4 1.1287n
L5 N4 N5 81.7578p
L6 N5 N6 57.5177p
R1 2 N1 2.4982
R2 2 N2 2.5011
R3 2 N3 1.3268
R4 2 N4 909.5526m
R5 2 N5 888.9213m
R6 2 N6 880.2481m
R7 2 N7 2.6427
R8 2 1 10g
.ends 
*******
.subckt 0402_744901051_5.1n 1 2
C1 1 N7 155.3952f
L1 1 N1 4.85n
L2 N1 N2 321.2646p
L3 N2 N3 96.3896p
L4 N3 N4 929.4816p
L5 N4 N5 85.5758p
L6 N5 N6 58.5814p
R1 2 N1 2.3968
R2 2 N2 1.6772
R3 2 N3 1.6304
R4 2 N4 1.2293
R5 2 N5 1.2078
R6 2 N6 1.1779
R7 2 N7 2.5604
R8 2 1 10g
.ends 
*******
.subckt 0402_744901056_5.6n 1 2
C1 1 N7 173.4310f
L1 1 N1 5.4n
L2 N1 N2 381.7743p
L3 N2 N3 114.8911p
L4 N3 N4 1.9707n
L5 N4 N5 85.6296p
L6 N5 N6 58.6080p
R1 2 N1 2.4123
R2 2 N2 1.6873
R3 2 N3 1.64
R4 2 N4 1.2271
R5 2 N5 1.2052
R6 2 N6 1.175
R7 2 N7 2.5606
R8 2 1 10g
.ends 
*******
.subckt 0402_744901058_5.8n 1 2
C1 1 N7 121.3f
L1 1 N1 5.5n
L2 N1 N2 338.3483p
L3 N2 N3 114.8422p
L4 N3 N4 1.9705n
L5 N4 N5 85.6284p
L6 N5 N6 58.6075p
R1 2 N1 2.4011
R2 2 N2 1.6863
R3 2 N3 1.6401
R4 2 N4 1.2272
R5 2 N5 1.2053
R6 2 N6 1.1751
R7 2 N7 2.5598
R8 2 1 10g
.ends 
*******
.subckt 0402_744901062_6.2n 1 2
C1 1 N7 113.487f
L1 1 N1 5.85n
L2 N1 N2 317.7346p
L3 N2 N3 113.7882p
L4 N3 N4 1.8645n
L5 N4 N5 85.1895p
L6 N5 N6 58.5004p
R1 2 N1 2.3308
R2 2 N2 1.5434
R3 2 N3 1.4774
R4 2 N4 1.2443
R5 2 N5 1.2264
R6 2 N6 1.1984
R7 2 N7 2.5615
R8 2 1 10g
.ends 
*******
.subckt 0402_744901068_6.8n 1 2
C1 1 N7 103.47f
L1 1 N1 6.42n
L2 N1 N2 430.2608p
L3 N2 N3 113.9423p
L4 N3 N4 1.8647n
L5 N4 N5 85.1923p
L6 N5 N6 58.5037p
R1 2 N1 3.3435
R2 2 N2 2.5599
R3 2 N3 1.5842
R4 2 N4 1.2486
R5 2 N5 1.2308
R6 2 N6 1.203
R7 2 N7 2.7604
R8 2 1 10g
.ends 
*******
.subckt 0402_744901072_7.2n 1 2
C1 1 N7 241.6367f
L1 1 N1 7n
L2 N1 N2 909.0220p
L3 N2 N3 3.4482n
L4 N3 N4 6.1424n
L5 N4 N5 121.9551p
L6 N5 N6 75.6623p
R1 2 N1 1.6929
R2 2 N2 1.3342
R3 2 N3 1.2721
R4 2 N4 2.4555
R5 2 N5 520.2094m
R6 2 N6 518.7389m
R7 2 N7 1.2510
R8 2 1 10g
.ends 
*******
.subckt 0402_744901082_8.2n 1 2
C1 1 N7 102.12f
L1 1 N1 7.8n
L2 N1 N2 720.0971p
L3 N2 N3 115.2093p
L4 N3 N4 1.8680n
L5 N4 N5 85.2048p
L6 N5 N6 58.5097p
R1 2 N1 3.3646
R2 2 N2 2.5754
R3 2 N3 1.6091
R4 2 N4 1.2504
R5 2 N5 1.2326
R6 2 N6 1.2049
R7 2 N7 2.7596
R8 2 1 10g
.ends 
*******
.subckt 0402_744901091_9.1n 1 2
C1 1 N7 195.2025f
L1 1 N1 8.3n
L2 N1 N2 595.9792p
L3 N2 N3 170.8678p
L4 N3 N4 1.8613n
L5 N4 N5 85.2322p
L6 N5 N6 58.5422p
R1 2 N1 3.3077
R2 2 N2 2.6003
R3 2 N3 1.6679
R4 2 N4 1.3266
R5 2 N5 1.3108
R6 2 N6 1.2864
R7 2 N7 2.7647
R8 2 1 10g
.ends 
*******
.subckt 0402_744901110_10n 1 2
C1 1 N7 134.2037f
L1 1 N1 9.3n
L2 N1 N2 628.2463p
L3 N2 N3 106.9797p
L4 N3 N4 2.0733n
L5 N4 N5 86.8456p
L6 N5 N6 58.9793p
R1 2 N1 6.2919
R2 2 N2 2.9291
R3 2 N3 4.7182
R4 2 N4 2.2176
R5 2 N5 2.2163
R6 2 N6 2.2094
R7 2 N7 5.4876
R8 2 1 10g
.ends 
*******
.subckt 0402_744901112_12n 1 2
C1 1 N7 153.1201f
L1 1 N1 11n
L2 N1 N2 791.3544p
L3 N2 N3 110.1428p
L4 N3 N4 2.3124n
L5 N4 N5 87.9496p
L6 N5 N6 59.2751p
R1 2 N1 6.287
R2 2 N2 3.0829
R3 2 N3 4.779
R4 2 N4 2.3463
R5 2 N5 2.3411
R6 2 N6 2.3336
R7 2 N7 5.4898
R8 2 1 10g
.ends 
*******
.subckt 0402_744901115_15n 1 2
C1 1 N7 320f
L1 1 N1 13.5n
L2 N1 N2 1.0748n
L3 N2 N3 110.8879p
L4 N3 N4 2.3303n
L5 N4 N5 88.0273p
L6 N5 N6 59.2910p
R1 2 N1 6.3115
R2 2 N2 3.1073
R3 2 N3 4.7872
R4 2 N4 2.3517
R5 2 N5 2.3463
R6 2 N6 2.3387
R7 2 N7 5.5093
R8 2 1 10g
.ends 
*******
.subckt 0402_744901118_18n 1 2
C1 1 N7 155.5383f
L1 1 N1 16n
L2 N1 N2 1.1981n
L3 N2 N3 298.0258p
L4 N3 N4 6.6345n
L5 N4 N5 355.9034p
L6 N5 N6 67.1343p
R1 2 N1 9.8409
R2 2 N2 5.8693
R3 2 N3 7.6285
R4 2 N4 5.6692
R5 2 N5 3.6435
R6 2 N6 3.6369
R7 2 N7 18.4088
R8 2 1 10g
.ends 
*******
.subckt 0402_744901122_22n 1 2
C1 1 N7 149.0896f
L1 1 N1 18n
L2 N1 N2 1.3676n
L3 N2 N3 298.6902p
L4 N3 N4 6.6313n
L5 N4 N5 355.8667p
L6 N5 N6 67.1344p
R1 2 N1 9.8557
R2 2 N2 5.8698
R3 2 N3 7.6288
R4 2 N4 5.6691
R5 2 N5 3.6433
R6 2 N6 3.6367
R7 2 N7 18.4083
R8 2 1 10g
.ends 
*******
.subckt 0402_744901127_27n 1 2
C1 1 N7 482.1453f
L1 1 N1 26.1n
L2 N1 N2 3.6452n
L3 N2 N3 5.8270n
L4 N3 N4 26.6208n
L5 N4 N5 100.7301p
L6 N5 N6 74.1350p
R1 2 N1 5.6776
R2 2 N2 2.0230
R3 2 N3 2.8378
R4 2 N4 3.9435
R5 2 N5 3.7842
R6 2 N6 3.7823
R7 2 N7 4.6763
R8 2 1 10g
.ends 
*******
