**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  SMT Power Inductor
* Matchcode:              WE-PD
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/27/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1030_7447713015_1.5u 1 2
Rp 1 2 672.674
Cp 1 2 3.599p
Rs 1 N3 0.0137
L1 N3 2 1.411u
.ends 1030_7447713015_1.5u
*******
.subckt 1030_7447713022_2.2u 1 2
Rp 1 2 945.477
Cp 1 2 2.803p
Rs 1 N3 0.0168
L1 N3 2 2.074u
.ends 1030_7447713022_2.2u
*******
.subckt 1030_7447713033_3.3u 1 2
Rp 1 2 1251
Cp 1 2 3.775p
Rs 1 N3 0.0204
L1 N3 2 3.005u
.ends 1030_7447713033_3.3u
*******
.subckt 1030_7447713047_4.7u 1 2
Rp 1 2 1701
Cp 1 2 4.595p
Rs 1 N3 0.026
L1 N3 2 4.271u
.ends 1030_7447713047_4.7u
*******
.subckt 1030_7447713082_8.2u 1 2
Rp 1 2 3617
Cp 1 2 4.502p
Rs 1 N3 0.041
L1 N3 2 7.276u
.ends 1030_7447713082_8.2u
*******
.subckt 1030_7447713100_10u 1 2
Rp 1 2 3554
Cp 1 2 4.934p
Rs 1 N3 0.0515
L1 N3 2 9.513u
.ends 1030_7447713100_10u
*******
.subckt 1030_7447713150_15u 1 2
Rp 1 2 5482
Cp 1 2 5.206p
Rs 1 N3 0.074
L1 N3 2 14.23u
.ends 1030_7447713150_15u
*******
.subckt 1030_7447713220_22u 1 2
Rp 1 2 8834
Cp 1 2 4.433p
Rs 1 N3 0.111
L1 N3 2 22.176u
.ends 1030_7447713220_22u
*******
.subckt 1030_7447713330_33u 1 2
Rp 1 2 12173
Cp 1 2 5.094p
Rs 1 N3 0.17
L1 N3 2 33.747u
.ends 1030_7447713330_33u
*******
.subckt 1030_7447713470_47u 1 2
Rp 1 2 13604
Cp 1 2 5.295p
Rs 1 N3 0.207
L1 N3 2 44.871u
.ends 1030_7447713470_47u
*******
.subckt 1030_7447713680_68u 1 2
Rp 1 2 19479
Cp 1 2 5.574p
Rs 1 N3 0.275
L1 N3 2 62.353u
.ends 1030_7447713680_68u
*******
.subckt 1030_7447713820_82u 1 2
Rp 1 2 25005
Cp 1 2 4.979p
Rs 1 N3 0.349
L1 N3 2 77.094u
.ends 1030_7447713820_82u
*******
.subckt 1030_7447713101_100u 1 2
Rp 1 2 30774
Cp 1 2 5.57p
Rs 1 N3 0.398
L1 N3 2 90.236u
.ends 1030_7447713101_100u
*******
.subckt 1030_7447713121_120u 1 2
Rp 1 2 40013
Cp 1 2 6.019p
Rs 1 N3 0.498
L1 N3 2 108.186u
.ends 1030_7447713121_120u
*******
.subckt 1030_7447713151_150u 1 2
Rp 1 2 46224
Cp 1 2 6.026p
Rs 1 N3 0.57
L1 N3 2 131.081u
.ends 1030_7447713151_150u
*******
.subckt 1030_7447713331_330u 1 2
Rp 1 2 72960
Cp 1 2 6.929p
Rs 1 N3 1.23
L1 N3 2 300.245u
.ends 1030_7447713331_330u
*******
.subckt 1030_7447713471_470u 1 2
Rp 1 2 88623
Cp 1 2 7.58p
Rs 1 N3 1.85
L1 N3 2 453.905u
.ends 1030_7447713471_470u
*******
.subckt 1030_7447713102_1000u 1 2
Rp 1 2 121895
Cp 1 2 8.544p
Rs 1 N3 4
L1 N3 2 957.63u
.ends 1030_7447713102_1000u
*******
.subckt 1050_7447714015_1.5u 1 2
Rp 1 2 696.48
Cp 1 2 3.69p
Rs 1 N3 0.00555
L1 N3 2 1.319u
.ends 1050_7447714015_1.5u
*******
.subckt 1050_7447714022_2.2u 1 2
Rp 1 2 1088
Cp 1 2 4.313p
Rs 1 N3 0.0068
L1 N3 2 2.019u
.ends 1050_7447714022_2.2u
*******
.subckt 1050_7447714033_3.3u 1 2
Rp 1 2 1748
Cp 1 2 4.94p
Rs 1 N3 0.0089
L1 N3 2 2.946u
.ends 1050_7447714033_3.3u
*******
.subckt 1050_7447714047_4.7u 1 2
Rp 1 2 2469
Cp 1 2 6.027p
Rs 1 N3 0.0104
L1 N3 2 4.148u
.ends 1050_7447714047_4.7u
*******
.subckt 1050_7447714056_5.6u 1 2
Rp 1 2 3639
Cp 1 2 6.084p
Rs 1 N3 0.012
L1 N3 2 5.401u
.ends 1050_7447714056_5.6u
*******
.subckt 1050_7447714068_6.8u 1 2
Rp 1 2 4349
Cp 1 2 7.2p
Rs 1 N3 0.0185
L1 N3 2 6.801u
.ends 1050_7447714068_6.8u
*******
.subckt 1050_7447714100_10u 1 2
Rp 1 2 6553
Cp 1 2 5.759p
Rs 1 N3 0.023
L1 N3 2 10.478u
.ends 1050_7447714100_10u
*******
.subckt 1050_7447714150_15u 1 2
Rp 1 2 9843
Cp 1 2 7.012p
Rs 1 N3 0.036
L1 N3 2 14.644u
.ends 1050_7447714150_15u
*******
.subckt 1050_7447714220_22u 1 2
Rp 1 2 12907
Cp 1 2 8.49p
Rs 1 N3 0.042
L1 N3 2 19.015u
.ends 1050_7447714220_22u
*******
.subckt 1050_7447714270_27u 1 2
Rp 1 2 16222
Cp 1 2 5.184p
Rs 1 N3 0.063
L1 N3 2 25.048u
.ends 1050_7447714270_27u
*******
.subckt 1050_7447714330_33u 1 2
Rp 1 2 18157
Cp 1 2 6.736p
Rs 1 N3 0.066
L1 N3 2 30.715u
.ends 1050_7447714330_33u
*******
.subckt 1050_7447714470_47u 1 2
Rp 1 2 25556
Cp 1 2 7.453p
Rs 1 N3 0.0825
L1 N3 2 45.428u
.ends 1050_7447714470_47u
*******
.subckt 1050_7447714560_56u 1 2
Rp 1 2 25720
Cp 1 2 6.476p
Rs 1 N3 0.101
L1 N3 2 52.405u
.ends 1050_7447714560_56u
*******
.subckt 1050_7447714680_68u 1 2
Rp 1 2 32590
Cp 1 2 6.803p
Rs 1 N3 0.11
L1 N3 2 61.871u
.ends 1050_7447714680_68u
*******
.subckt 1050_7447714820_82u 1 2
Rp 1 2 33435
Cp 1 2 7.917p
Rs 1 N3 0.147
L1 N3 2 78.213u
.ends 1050_7447714820_82u
*******
.subckt 1050_7447714101_100u 1 2
Rp 1 2 33721
Cp 1 2 8.231p
Rs 1 N3 0.165
L1 N3 2 93.461u
.ends 1050_7447714101_100u
*******
.subckt 1050_7447714151_150u 1 2
Rp 1 2 53063
Cp 1 2 9.967p
Rs 1 N3 0.251
L1 N3 2 138.62u
.ends 1050_7447714151_150u
*******
.subckt 1050_7447714221_220u 1 2
Rp 1 2 61488
Cp 1 2 6.439p
Rs 1 N3 0.366
L1 N3 2 196.516u
.ends 1050_7447714221_220u
*******
.subckt 1050_7447714331_330u 1 2
Rp 1 2 79107
Cp 1 2 9.655p
Rs 1 N3 0.655
L1 N3 2 325.418u
.ends 1050_7447714331_330u
*******
.subckt 1050_7447714471_470u 1 2
Rp 1 2 77358
Cp 1 2 10.702p
Rs 1 N3 0.96
L1 N3 2 441.117u
.ends 1050_7447714471_470u
*******
.subckt 1050_7447714681_680u 1 2
Rp 1 2 92097
Cp 1 2 11.336p
Rs 1 N3 1.22
L1 N3 2 631.718u
.ends 1050_7447714681_680u
*******
.subckt 1050_7447714102_1000u 1 2
Rp 1 2 180643
Cp 1 2 7.59p
Rs 1 N3 1.86
L1 N3 2 908.799u
.ends 1050_7447714102_1000u
*******
.subckt 1050P_7447714152_1500u 1 2
Rp 1 2 281646
Cp 1 2 11.328p
Rs 1 N3 3.04
L1 N3 2 1431u
.ends 1050P_7447714152_1500u
*******
.subckt 1210_7447709001_1u 1 2
Rp 1 2 2176.6207769
Cp 1 2 2.24744833282p
Rs 1 N3 0.004
L1 N3 2 0.888311902286u
.ends 1210_7447709001_1u
*******
.subckt 1210_7447709002_2.2u 1 2
Rp 1 2 4137.02857985
Cp 1 2 2.99089969563p
Rs 1 N3 0.005
L1 N3 2 2.04316893219u
.ends 1210_7447709002_2.2u
*******
.subckt 1210_7447709003_3.5u 1 2
Rp 1 2 4975.69579666
Cp 1 2 4.15650993146p
Rs 1 N3 0.006
L1 N3 2 3.04371144857u
.ends 1210_7447709003_3.5u
*******
.subckt 1210_7447709004_4.7u 1 2
Rp 1 2 5047
Cp 1 2 6.87p
Rs 1 N3 0.007
L1 N3 2 3.84u
.ends 1210_7447709004_4.7u
*******
.subckt 1210_7447709006_6.8u 1 2
Rp 1 2 8250.62950059
Cp 1 2 7.73395856798p
Rs 1 N3 0.009
L1 N3 2 6.30631538292u
.ends 1210_7447709006_6.8u
*******
.subckt 1210_7447709100_10u 1 2
Rp 1 2 11546.6960325
Cp 1 2 7.27315529525p
Rs 1 N3 0.013
L1 N3 2 9.52800542568u
.ends 1210_7447709100_10u
*******
.subckt 1210_7447709150_15u 1 2
Rp 1 2 15765.1384684
Cp 1 2 7.13382716865p
Rs 1 N3 0.021
L1 N3 2 12.6985405468u
.ends 1210_7447709150_15u
*******
.subckt 1210_7447709220_22u 1 2
Rp 1 2 13263
Cp 1 2 14.26p
Rs 1 N3 0.023
L1 N3 2 18.65u
.ends 1210_7447709220_22u
*******
.subckt 1210_7447709270_27u 1 2
Rp 1 2 29129.0712954
Cp 1 2 13.9416435215p
Rs 1 N3 0.03
L1 N3 2 23.0051014632u
.ends 1210_7447709270_27u
*******
.subckt 1210_7447709330_33u 1 2
Rp 1 2 30639.6783453
Cp 1 2 13.0681350616p
Rs 1 N3 0.037
L1 N3 2 31.196u
.ends 1210_7447709330_33u
*******
.subckt 1210_7447709390_39u 1 2
Rp 1 2 36480.6887288
Cp 1 2 16.6752475935p
Rs 1 N3 0.044
L1 N3 2 31.879u
.ends 1210_7447709390_39u
*******
.subckt 1210_7447709470_47u 1 2
Rp 1 2 43179.7160489
Cp 1 2 15.5579429534p
Rs 1 N3 0.046
L1 N3 2 44.953u
.ends 1210_7447709470_47u
*******
.subckt 1210_7447709680_68u 1 2
Rp 1 2 65987.2147297
Cp 1 2 15.6960659854p
Rs 1 N3 0.069
L1 N3 2 55.0105245384u
.ends 1210_7447709680_68u
*******
.subckt 1210_7447709820_82u 1 2
Rp 1 2 39761
Cp 1 2 15.516p
Rs 1 N3 0.0905
L1 N3 2 79.63u
.ends 1210_7447709820_82u
*******
.subckt 1210_7447709101_100u 1 2
Rp 1 2 59146
Cp 1 2 18.224p
Rs 1 N3 0.1
L1 N3 2 93.766u
.ends 1210_7447709101_100u
*******
.subckt 1210_7447709151_150u 1 2
Rp 1 2 82598.270635
Cp 1 2 14.2781138855p
Rs 1 N3 0.151
L1 N3 2 144.009u
.ends 1210_7447709151_150u
*******
.subckt 1210_7447709221_220u 1 2
Rp 1 2 91179.4137734
Cp 1 2 16.3697778895p
Rs 1 N3 0.193
L1 N3 2 212.529u
.ends 1210_7447709221_220u
*******
.subckt 1210_7447709271_270u 1 2
Rp 1 2 99265.0050729
Cp 1 2 18.0619283051p
Rs 1 N3 0.248
L1 N3 2 256u
.ends 1210_7447709271_270u
*******
.subckt 1210_7447709331_330u 1 2
Rp 1 2 90525.0521166
Cp 1 2 20.1460207887p
Rs 1 N3 0.363
L1 N3 2 327.159u
.ends 1210_7447709331_330u
*******
.subckt 1210_7447709471_470u 1 2
Rp 1 2 105258.807914
Cp 1 2 20.5928638778p
Rs 1 N3 0.437
L1 N3 2 436.648u
.ends 1210_7447709471_470u
*******
.subckt 1210_7447709681_680u 1 2
Rp 1 2 120411.679361
Cp 1 2 19.3385293438p
Rs 1 N3 0.66
L1 N3 2 668.961u
.ends 1210_7447709681_680u
*******
.subckt 1210_7447709821_820u 1 2
Rp 1 2 117117.877304
Cp 1 2 21.7929604862p
Rs 1 N3 0.815
L1 N3 2 799.794u
.ends 1210_7447709821_820u
*******
.subckt 1210_7447709102_1000u 1 2
Rp 1 2 103052
Cp 1 2 21.42p
Rs 1 N3 0.93
L1 N3 2 982.946u
.ends 1210_7447709102_1000u
*******
.subckt 1210_7447709152_1500u 1 2
Rp 1 2 171070
Cp 1 2 25.56p
Rs 1 N3 1.8
L1 N3 2 1423u
.ends 1210_7447709152_1500u
*******
.subckt 1210_7447709222_2200u 1 2
Rp 1 2 200000
Cp 1 2 30p
Rs 1 N3 3.25
L1 N3 2 2122u
.ends 1210_7447709222_2200u
*******
.subckt 1245_7447715906_0.6u 1 2
Rp 1 2 1308.28965673
Cp 1 2 2.223341372p
Rs 1 N3 0.0045
L1 N3 2 0.464397869128u
.ends 1245_7447715906_0.6u
*******
.subckt 1245_7447715910_1u 1 2
Rp 1 2 2427.45429051
Cp 1 2 3.07393402306p
Rs 1 N3 0.0055
L1 N3 2 0.874032032284u
.ends 1245_7447715910_1u
*******
.subckt 1245_7447715001_1.8u 1 2
Rp 1 2 3556.81358598
Cp 1 2 3.49530401983p
Rs 1 N3 0.0075
L1 N3 2 1.5713563659u
.ends 1245_7447715001_1.8u
*******
.subckt 1245_7447715002_2.5u 1 2
Rp 1 2 3968.08010791
Cp 1 2 3.66763216981p
Rs 1 N3 0.0085
L1 N3 2 2.51732267391u
.ends 1245_7447715002_2.5u
*******
.subckt 1245_7447715003_3.3u 1 2
Rp 1 2 6578.47426969
Cp 1 2 4.39654551772p
Rs 1 N3 0.0115
L1 N3 2 2.88851569677u
.ends 1245_7447715003_3.3u
*******
.subckt 1245_7447715004_4.7u 1 2
Rp 1 2 8219.38035441
Cp 1 2 4.06523390514p
Rs 1 N3 0.0135
L1 N3 2 3.75692461883u
.ends 1245_7447715004_4.7u
*******
.subckt 1245_7447715006_6.8u 1 2
Rp 1 2 11078.5420015
Cp 1 2 4.29910927901p
Rs 1 N3 0.02
L1 N3 2 6.87526199363u
.ends 1245_7447715006_6.8u
*******
.subckt 1245_7447715100_10u 1 2
Rp 1 2 15515.0080042
Cp 1 2 4.83057400324p
Rs 1 N3 0.025
L1 N3 2 9.01972200031u
.ends 1245_7447715100_10u
*******
.subckt 1245_7447715120_12u 1 2
Rp 1 2 16500.8527686
Cp 1 2 4.85170401496p
Rs 1 N3 0.03
L1 N3 2 10.705444972u
.ends 1245_7447715120_12u
*******
.subckt 1245_7447715180_18u 1 2
Rp 1 2 20313.2567777
Cp 1 2 5.45940158137p
Rs 1 N3 0.037
L1 N3 2 13.0855292701u
.ends 1245_7447715180_18u
*******
.subckt 1245_7447715220_22u 1 2
Rp 1 2 26167.9513606
Cp 1 2 5.27045194002p
Rs 1 N3 0.045
L1 N3 2 17.3598966267u
.ends 1245_7447715220_22u
*******
.subckt 1245_7447715330_33u 1 2
Rp 1 2 35410.3838309
Cp 1 2 5.06743999531p
Rs 1 N3 0.075
L1 N3 2 25.7301392598u
.ends 1245_7447715330_33u
*******
.subckt 1245_7447715470_47u 1 2
Rp 1 2 52874.4211867
Cp 1 2 5.23820249993p
Rs 1 N3 0.105
L1 N3 2 37.929937389u
.ends 1245_7447715470_47u
*******
.subckt 1245_7447715101_100u 1 2
Rp 1 2 96148.7175854
Cp 1 2 5.79622090066p
Rs 1 N3 0.25
L1 N3 2 80.390308916u
.ends 1245_7447715101_100u
*******
.subckt 1245_7447715221_220u 1 2
Rp 1 2 130584.615405
Cp 1 2 5.82141733606p
Rs 1 N3 0.46
L1 N3 2 167.025850479u
.ends 1245_7447715221_220u
*******
.subckt 1260_744771010_1u 1 2
Rp 1 2 1862
Cp 1 2 3.48p
Rs 1 N3 0.003
L1 N3 2 0.889329u
.ends 1260_744771010_1u
*******
.subckt 1260_7447706015_1.5u 1 2
Rp 1 2 665
Cp 1 2 7.3p
Rs 1 N3 0.005
L1 N3 2 1.363u
.ends 1260_7447706015_1.5u
*******
.subckt 1260_744771001_1.5u 1 2
Rp 1 2 2665
Cp 1 2 4.377p
Rs 1 N3 0.004
L1 N3 2 1.402u
.ends 1260_744771001_1.5u
*******
.subckt 1260_744771002_2.2u 1 2
Rp 1 2 3696
Cp 1 2 4.203p
Rs 1 N3 0.005
L1 N3 2 2.069u
.ends 1260_744771002_2.2u
*******
.subckt 1260_7447706022_2.2u 1 2
Rp 1 2 1109
Cp 1 2 6.96p
Rs 1 N3 0.0062
L1 N3 2 2.251u
.ends 1260_7447706022_2.2u
*******
.subckt 1260_744771003_3.5u 1 2
Rp 1 2 4638
Cp 1 2 5.297p
Rs 1 N3 0.0055
L1 N3 2 2.724u
.ends 1260_744771003_3.5u
*******
.subckt 1260_7447706033_3.3u 1 2
Rp 1 2 1721
Cp 1 2 7.452p
Rs 1 N3 0.0075
L1 N3 2 3.28u
.ends 1260_7447706033_3.3u
*******
.subckt 1260_744771004_4.7u 1 2
Rp 1 2 5213
Cp 1 2 5.126p
Rs 1 N3 0.0085
L1 N3 2 3.746u
.ends 1260_744771004_4.7u
*******
.subckt 1260_7447706047_4.7u 1 2
Rp 1 2 2353
Cp 1 2 7.333p
Rs 1 N3 0.009
L1 N3 2 4.594u
.ends 1260_7447706047_4.7u
*******
.subckt 1260_7447706062_6.2u 1 2
Rp 1 2 3316
Cp 1 2 8.206p
Rs 1 N3 0.012
L1 N3 2 6.122u
.ends 1260_7447706062_6.2u
*******
.subckt 1260_744771008_8.2u 1 2
Rp 1 2 9391
Cp 1 2 5.647p
Rs 1 N3 0.0155
L1 N3 2 6.458u
.ends 1260_744771008_8.2u
*******
.subckt 1260_744771006_6.8u 1 2
Rp 1 2 8031
Cp 1 2 5.64p
Rs 1 N3 0.014
L1 N3 2 6.463u
.ends 1260_744771006_6.8u
*******
.subckt 1260_7447706100_10u 1 2
Rp 1 2 5174
Cp 1 2 8.558p
Rs 1 N3 0.0163
L1 N3 2 9.54u
.ends 1260_7447706100_10u
*******
.subckt 1260_74477110_10u 1 2
Rp 1 2 11359
Cp 1 2 5.93p
Rs 1 N3 0.0185
L1 N3 2 9.753u
.ends 1260_74477110_10u
*******
.subckt 1260_744771112_12u 1 2
Rp 1 2 13114
Cp 1 2 6.319p
Rs 1 N3 0.02
L1 N3 2 11.334u
.ends 1260_744771112_12u
*******
.subckt 1260_744771115_15u 1 2
Rp 1 2 13381
Cp 1 2 6.382p
Rs 1 N3 0.022
L1 N3 2 12.996u
.ends 1260_744771115_15u
*******
.subckt 1260_7447706150_15u 1 2
Rp 1 2 7898
Cp 1 2 9.234p
Rs 1 N3 0.0229
L1 N3 2 14.117u
.ends 1260_7447706150_15u
*******
.subckt 1260_744771118_18u 1 2
Rp 1 2 14024
Cp 1 2 5.88p
Rs 1 N3 0.024
L1 N3 2 14.994u
.ends 1260_744771118_18u
*******
.subckt 1260_744771122_22u 1 2
Rp 1 2 17438
Cp 1 2 6.037p
Rs 1 N3 0.03
L1 N3 2 18.295u
.ends 1260_744771122_22u
*******
.subckt 1260_7447706220_22u 1 2
Rp 1 2 11306
Cp 1 2 9.325p
Rs 1 N3 0.0343
L1 N3 2 22.406u
.ends 1260_7447706220_22u
*******
.subckt 1260_744771127_27u 1 2
Rp 1 2 19869
Cp 1 2 6.308p
Rs 1 N3 0.037
L1 N3 2 23.729u
.ends 1260_744771127_27u
*******
.subckt 1260_744771133_33u 1 2
Rp 1 2 19960
Cp 1 2 6.391p
Rs 1 N3 0.049
L1 N3 2 30.263u
.ends 1260_744771133_33u
*******
.subckt 1260_7447706330_33u 1 2
Rp 1 2 14360
Cp 1 2 9.175p
Rs 1 N3 0.0508
L1 N3 2 32.823u
.ends 1260_7447706330_33u
*******
.subckt 1260_744771139_39u 1 2
Rp 1 2 23972
Cp 1 2 6.972p
Rs 1 N3 0.057
L1 N3 2 35.479u
.ends 1260_744771139_39u
*******
.subckt 1260_744771147_47u 1 2
Rp 1 2 26156
Cp 1 2 6.858p
Rs 1 N3 0.064
L1 N3 2 39.609u
.ends 1260_744771147_47u
*******
.subckt 1260_7447706470_47u 1 2
Rp 1 2 19493
Cp 1 2 10.085p
Rs 1 N3 0.0612
L1 N3 2 44.161u
.ends 1260_7447706470_47u
*******
.subckt 1260_744771156_56u 1 2
Rp 1 2 35043
Cp 1 2 6.797p
Rs 1 N3 0.077
L1 N3 2 51.171u
.ends 1260_744771156_56u
*******
.subckt 1260_744771168_68u 1 2
Rp 1 2 38057
Cp 1 2 7.521p
Rs 1 N3 0.086
L1 N3 2 60.094u
.ends 1260_744771168_68u
*******
.subckt 1260_7447706680_68u 1 2
Rp 1 2 25360
Cp 1 2 9.53p
Rs 1 N3 0.082
L1 N3 2 64.035u
.ends 1260_7447706680_68u
*******
.subckt 1260_744771182_82u 1 2
Rp 1 2 47497
Cp 1 2 7.093p
Rs 1 N3 0.112
L1 N3 2 75.648u
.ends 1260_744771182_82u
*******
.subckt 1260_74477120_100u 1 2
Rp 1 2 52186
Cp 1 2 7.386p
Rs 1 N3 0.135
L1 N3 2 90.601u
.ends 1260_74477120_100u
*******
.subckt 1260_7447706101_100u 1 2
Rp 1 2 34132
Cp 1 2 10.21p
Rs 1 N3 0.122
L1 N3 2 90.851u
.ends 1260_7447706101_100u
*******
.subckt 1260_744771212_120u 1 2
Rp 1 2 55504
Cp 1 2 6.865p
Rs 1 N3 0.15
L1 N3 2 108.278u
.ends 1260_744771212_120u
*******
.subckt 1260_744771215_150u 1 2
Rp 1 2 68654
Cp 1 2 7.441p
Rs 1 N3 0.185
L1 N3 2 135.504u
.ends 1260_744771215_150u
*******
.subckt 1260_7447706151_150u 1 2
Rp 1 2 43015
Cp 1 2 10.304p
Rs 1 N3 0.175
L1 N3 2 138.623u
.ends 1260_7447706151_150u
*******
.subckt 1260_744771218_180u 1 2
Rp 1 2 75000
Cp 1 2 7.649p
Rs 1 N3 0.23
L1 N3 2 156.586u
.ends 1260_744771218_180u
*******
.subckt 1260_744771220_220u 1 2
Rp 1 2 77433
Cp 1 2 7.283p
Rs 1 N3 0.28
L1 N3 2 202.464u
.ends 1260_744771220_220u
*******
.subckt 1260_7447706221_220u 1 2
Rp 1 2 61324
Cp 1 2 11.14p
Rs 1 N3 0.273
L1 N3 2 206.417u
.ends 1260_7447706221_220u
*******
.subckt 1260_744771270_270u 1 2
Rp 1 2 80000
Cp 1 2 7.5p
Rs 1 N3 0.33
L1 N3 2 246.708u
.ends 1260_744771270_270u
*******
.subckt 1260_744771233_330u 1 2
Rp 1 2 93949
Cp 1 2 7.976p
Rs 1 N3 0.41
L1 N3 2 300.162u
.ends 1260_744771233_330u
*******
.subckt 1260_7447706331_330u 1 2
Rp 1 2 77487
Cp 1 2 11.608p
Rs 1 N3 0.395
L1 N3 2 313.836u
.ends 1260_7447706331_330u
*******
.subckt 1260_744771239_390u 1 2
Rp 1 2 96846
Cp 1 2 8.1p
Rs 1 N3 0.54
L1 N3 2 360.487u
.ends 1260_744771239_390u
*******
.subckt 1260_74477124_470u 1 2
Rp 1 2 121785
Cp 1 2 7.901p
Rs 1 N3 0.59
L1 N3 2 431.521u
.ends 1260_74477124_470u
*******
.subckt 1260_7447706471_470u 1 2
Rp 1 2 79506
Cp 1 2 11.059p
Rs 1 N3 0.543
L1 N3 2 445.248u
.ends 1260_7447706471_470u
*******
.subckt 1260_74477125_560u 1 2
Rp 1 2 124884
Cp 1 2 7.961p
Rs 1 N3 0.74
L1 N3 2 530.155u
.ends 1260_74477125_560u
*******
.subckt 1260_74477126_680u 1 2
Rp 1 2 136460
Cp 1 2 7.095p
Rs 1 N3 0.85
L1 N3 2 632.579u
.ends 1260_74477126_680u
*******
.subckt 1260_7447706681_680u 1 2
Rp 1 2 103448
Cp 1 2 12.098p
Rs 1 N3 0.78
L1 N3 2 657.541u
.ends 1260_7447706681_680u
*******
.subckt 1260_74477128_820u 1 2
Rp 1 2 139306
Cp 1 2 7.059p
Rs 1 N3 0.98
L1 N3 2 764.395u
.ends 1260_74477128_820u
*******
.subckt 1260_7447706102_1000u 1 2
Rp 1 2 118912
Cp 1 2 12.776p
Rs 1 N3 1.15
L1 N3 2 943.548u
.ends 1260_7447706102_1000u
*******
.subckt 1260_74477130_1000u 1 2
Rp 1 2 176070
Cp 1 2 8.008p
Rs 1 N3 1.33
L1 N3 2 961u
.ends 1260_74477130_1000u
*******
.subckt 1280_74477009_0.47u 1 2
Rp 1 2 1045
Cp 1 2 4.301p
Rs 1 N3 0.0017
L1 N3 2 0.426471u
.ends 1280_74477009_0.47u
*******
.subckt 1280_74477008_0.75u 1 2
Rp 1 2 1844
Cp 1 2 2.903p
Rs 1 N3 0.0032
L1 N3 2 0.723257u
.ends 1280_74477008_0.75u
*******
.subckt 1280_74477001_1.2u 1 2
Rp 1 2 2329
Cp 1 2 13p
Rs 1 N3 0.0046
L1 N3 2 0.96686u
.ends 1280_74477001_1.2u
*******
.subckt 1280_744770015_1.5u 1 2
Rp 1 2 2509
Cp 1 2 11.5p
Rs 1 N3 0.0032
L1 N3 2 1.226u
.ends 1280_744770015_1.5u
*******
.subckt 1280_7447707015_1.5u 1 2
Rp 1 2 743
Cp 1 2 8.11p
Rs 1 N3 0.0046
L1 N3 2 1.289u
.ends 1280_7447707015_1.5u
*******
.subckt 1280_7447707022_2.2u 1 2
Rp 1 2 1218
Cp 1 2 6.996p
Rs 1 N3 0.0057
L1 N3 2 2.08u
.ends 1280_7447707022_2.2u
*******
.subckt 1280_74477002_2.4u 1 2
Rp 1 2 3879
Cp 1 2 7.08p
Rs 1 N3 0.0063
L1 N3 2 2.136u
.ends 1280_74477002_2.4u
*******
.subckt 1280_7447707033_3.3u 1 2
Rp 1 2 1847
Cp 1 2 7.991p
Rs 1 N3 0.0075
L1 N3 2 3.026u
.ends 1280_7447707033_3.3u
*******
.subckt 1280_74477003_3.5u 1 2
Rp 1 2 3620
Cp 1 2 4.974p
Rs 1 N3 0.008
L1 N3 2 3.814u
.ends 1280_74477003_3.5u
*******
.subckt 1280_7447707047_4.7u 1 2
Rp 1 2 2486
Cp 1 2 7.593p
Rs 1 N3 0.0085
L1 N3 2 4.012u
.ends 1280_7447707047_4.7u
*******
.subckt 1280_74477004_4.7u 1 2
Rp 1 2 7007
Cp 1 2 5.182p
Rs 1 N3 0.009
L1 N3 2 4.982u
.ends 1280_74477004_4.7u
*******
.subckt 1280_74477005_5.6u 1 2
Rp 1 2 5511
Cp 1 2 8p
Rs 1 N3 0.0105
L1 N3 2 5.464u
.ends 1280_74477005_5.6u
*******
.subckt 1280_74477006_6.1u 1 2
Rp 1 2 4617
Cp 1 2 6.759p
Rs 1 N3 0.011
L1 N3 2 6.063u
.ends 1280_74477006_6.1u
*******
.subckt 1280_74477007_7.6u 1 2
Rp 1 2 5744
Cp 1 2 8.653p
Rs 1 N3 0.0115
L1 N3 2 6.848u
.ends 1280_74477007_7.6u
*******
.subckt 1280_7447707068_6.8u 1 2
Rp 1 2 4411
Cp 1 2 9.915p
Rs 1 N3 0.0118
L1 N3 2 6.979u
.ends 1280_7447707068_6.8u
*******
.subckt 1280_74477010_10u 1 2
Rp 1 2 5267
Cp 1 2 8.638p
Rs 1 N3 0.015
L1 N3 2 8.785u
.ends 1280_74477010_10u
*******
.subckt 1280_7447707100_10u 1 2
Rp 1 2 6455
Cp 1 2 10.234p
Rs 1 N3 0.018
L1 N3 2 10.839u
.ends 1280_7447707100_10u
*******
.subckt 1280_744770112_12u 1 2
Rp 1 2 9991
Cp 1 2 8.834p
Rs 1 N3 0.016
L1 N3 2 11.559u
.ends 1280_744770112_12u
*******
.subckt 1280_744770115_15u 1 2
Rp 1 2 10951
Cp 1 2 10.107p
Rs 1 N3 0.018
L1 N3 2 12.42u
.ends 1280_744770115_15u
*******
.subckt 1280_7447707150_15u 1 2
Rp 1 2 8882
Cp 1 2 9.911p
Rs 1 N3 0.023
L1 N3 2 14.539u
.ends 1280_7447707150_15u
*******
.subckt 1280_744770118_18u 1 2
Rp 1 2 16340
Cp 1 2 8.407p
Rs 1 N3 0.025
L1 N3 2 17.889u
.ends 1280_744770118_18u
*******
.subckt 1280_7447707220_22u 1 2
Rp 1 2 12927
Cp 1 2 11.652p
Rs 1 N3 0.0315
L1 N3 2 20.747u
.ends 1280_7447707220_22u
*******
.subckt 1280_744770122_22u 1 2
Rp 1 2 19687
Cp 1 2 8.266p
Rs 1 N3 0.029
L1 N3 2 23.064u
.ends 1280_744770122_22u
*******
.subckt 1280_744770127_27u 1 2
Rp 1 2 16374
Cp 1 2 10.144p
Rs 1 N3 0.031
L1 N3 2 23.712u
.ends 1280_744770127_27u
*******
.subckt 1280_744770133_33u 1 2
Rp 1 2 17739
Cp 1 2 11.303p
Rs 1 N3 0.044
L1 N3 2 31.196u
.ends 1280_744770133_33u
*******
.subckt 1280_744770139_39u 1 2
Rp 1 2 22274
Cp 1 2 11.375p
Rs 1 N3 0.047
L1 N3 2 31.879u
.ends 1280_744770139_39u
*******
.subckt 1280_7447707330_33u 1 2
Rp 1 2 16036
Cp 1 2 11.112p
Rs 1 N3 0.0465
L1 N3 2 32.942u
.ends 1280_7447707330_33u
*******
.subckt 1280_7447707470_47u 1 2
Rp 1 2 21764
Cp 1 2 10.823p
Rs 1 N3 0.055
L1 N3 2 44.771u
.ends 1280_7447707470_47u
*******
.subckt 1280_744770147_47u 1 2
Rp 1 2 21959
Cp 1 2 9.148p
Rs 1 N3 0.053
L1 N3 2 44.953u
.ends 1280_744770147_47u
*******
.subckt 1280_744770156_56u 1 2
Rp 1 2 26781
Cp 1 2 9.998p
Rs 1 N3 0.059
L1 N3 2 50.957u
.ends 1280_744770156_56u
*******
.subckt 1280_744770168_68u 1 2
Rp 1 2 43066
Cp 1 2 10.899p
Rs 1 N3 0.076
L1 N3 2 61.924u
.ends 1280_744770168_68u
*******
.subckt 1280_7447707680_68u 1 2
Rp 1 2 26176
Cp 1 2 12.896p
Rs 1 N3 0.078
L1 N3 2 64.484u
.ends 1280_7447707680_68u
*******
.subckt 1280_744770182_82u 1 2
Rp 1 2 42188
Cp 1 2 24.9p
Rs 1 N3 0.086
L1 N3 2 79.63u
.ends 1280_744770182_82u
*******
.subckt 1280_74477020_100u 1 2
Rp 1 2 43243
Cp 1 2 9.795p
Rs 1 N3 0.117
L1 N3 2 93.766u
.ends 1280_74477020_100u
*******
.subckt 1280_7447707101_100u 1 2
Rp 1 2 46275
Cp 1 2 13.986p
Rs 1 N3 0.105
L1 N3 2 95.116u
.ends 1280_7447707101_100u
*******
.subckt 1280_7447707151_150u 1 2
Rp 1 2 52634
Cp 1 2 14.585p
Rs 1 N3 0.165
L1 N3 2 138.718u
.ends 1280_7447707151_150u
*******
.subckt 1280_744770215_150u 1 2
Rp 1 2 65343
Cp 1 2 19.585p
Rs 1 N3 0.145
L1 N3 2 144.009u
.ends 1280_744770215_150u
*******
.subckt 1280P_7447707181_180u 1 2
Rp 1 2 58634
Cp 1 2 14.785p
Rs 1 N3 0.225
L1 N3 2 168.718u
.ends 1280P_7447707181_180u
*******
.subckt 1280_744770218_180u 1 2
Rp 1 2 57579
Cp 1 2 8.108p
Rs 1 N3 0.182
L1 N3 2 179.242u
.ends 1280_744770218_180u
*******
.subckt 1280_7447707221_220u 1 2
Rp 1 2 61530
Cp 1 2 14.854p
Rs 1 N3 0.24
L1 N3 2 200.746u
.ends 1280_7447707221_220u
*******
.subckt 1280_744770222_220u 1 2
Rp 1 2 81630
Cp 1 2 8.317p
Rs 1 N3 0.23
L1 N3 2 212.529u
.ends 1280_744770222_220u
*******
.subckt 1280_7447707331_330u 1 2
Rp 1 2 73048
Cp 1 2 17.669p
Rs 1 N3 0.372
L1 N3 2 306.58u
.ends 1280_7447707331_330u
*******
.subckt 1280_744770233_330u 1 2
Rp 1 2 83993
Cp 1 2 8.56p
Rs 1 N3 0.345
L1 N3 2 327.159u
.ends 1280_744770233_330u
*******
.subckt 1280_744770247_470u 1 2
Rp 1 2 117817
Cp 1 2 8.535p
Rs 1 N3 0.45
L1 N3 2 436.648u
.ends 1280_744770247_470u
*******
.subckt 1280_7447707471_470u 1 2
Rp 1 2 87039
Cp 1 2 15.174p
Rs 1 N3 0.49
L1 N3 2 451.177u
.ends 1280_7447707471_470u
*******
.subckt 1280P_7447707561_560u 1 2
Rp 1 2 92000
Cp 1 2 15.2p
Rs 1 N3 0.58
L1 N3 2 527u
.ends 1280P_7447707561_560u
*******
.subckt 1280_744770256_560u 1 2
Rp 1 2 119841
Cp 1 2 7.43p
Rs 1 N3 0.57
L1 N3 2 546.802u
.ends 1280_744770256_560u
*******
.subckt 1280_7447707681_680u 1 2
Rp 1 2 96849
Cp 1 2 17.639p
Rs 1 N3 0.7
L1 N3 2 640.731u
.ends 1280_7447707681_680u
*******
.subckt 1280_744770268_680u 1 2
Rp 1 2 103542
Cp 1 2 7.85p
Rs 1 N3 0.78
L1 N3 2 668.961u
.ends 1280_744770268_680u
*******
.subckt 1280_744770282_820u 1 2
Rp 1 2 149541
Cp 1 2 8p
Rs 1 N3 0.87
L1 N3 2 799.794u
.ends 1280_744770282_820u
*******
.subckt 1280_7447707102_1000u 1 2
Rp 1 2 112243
Cp 1 2 17.971p
Rs 1 N3 0.985
L1 N3 2 952.938u
.ends 1280_7447707102_1000u
*******
.subckt 1280_74477030_1000u 1 2
Rp 1 2 145822
Cp 1 2 8.178p
Rs 1 N3 0.98
L1 N3 2 982.946u
.ends 1280_74477030_1000u
*******
.subckt 1510_7447704150_15u 1 2
Rp 1 2 11219
Cp 1 2 4.694p
Rs 1 N3 0.0195
L1 N3 2 12.92u
.ends 1510_7447704150_15u
*******
.subckt 1510_7447704220_22u 1 2
Rp 1 2 13326
Cp 1 2 9.74p
Rs 1 N3 0.025
L1 N3 2 19.837u
.ends 1510_7447704220_22u
*******
.subckt 1510_7447704471_470u 1 2
Rp 1 2 77780
Cp 1 2 20.119p
Rs 1 N3 0.425
L1 N3 2 420.593u
.ends 1510_7447704471_470u
*******
.subckt 6033_7447785001_1u 1 2
Rp 1 2 2216.77027065
Cp 1 2 0.857843400666p
Rs 1 N3 0.031
L1 N3 2 0.967255025011u
.ends 6033_7447785001_1u
*******
.subckt 6033_7447785002_2.2u 1 2
Rp 1 2 4378.30426868
Cp 1 2 1.81548178904p
Rs 1 N3 0.043
L1 N3 2 2.15314312624u
.ends 6033_7447785002_2.2u
*******
.subckt 6033_7447785003_3.3u 1 2
Rp 1 2 5378.14539148
Cp 1 2 2.0293197902p
Rs 1 N3 0.043
L1 N3 2 2.7563697661u
.ends 6033_7447785003_3.3u
*******
.subckt 6033_7447785004_4.7u 1 2
Rp 1 2 6419.16347886
Cp 1 2 2.18658481122p
Rs 1 N3 0.06
L1 N3 2 4.16756573005u
.ends 6033_7447785004_4.7u
*******
.subckt 6033_7447785006_6.8u 1 2
Rp 1 2 8506.21069778
Cp 1 2 2.12954534656p
Rs 1 N3 0.079
L1 N3 2 6.05071959927u
.ends 6033_7447785006_6.8u
*******
.subckt 6033_744778510_10u 1 2
Rp 1 2 12213.3283534
Cp 1 2 2.46060321425p
Rs 1 N3 0.1
L1 N3 2 8.79321625609u
.ends 6033_744778510_10u
*******
.subckt 6033_7447785115_15u 1 2
Rp 1 2 13553.342485
Cp 1 2 2.64078545593p
Rs 1 N3 0.165
L1 N3 2 14.7022745416u
.ends 6033_7447785115_15u
*******
.subckt 6033_7447785122_22u 1 2
Rp 1 2 21477.817611
Cp 1 2 2.33541671451p
Rs 1 N3 0.21
L1 N3 2 19.4251211974u
.ends 6033_7447785122_22u
*******
.subckt 6033_7447785127_27u 1 2
Rp 1 2 18720
Cp 1 2 2.76p
Rs 1 N3 0.3
L1 N3 2 25.123u
.ends 6033_7447785127_27u
*******
.subckt 6033_7447785133_33u 1 2
Rp 1 2 24630
Cp 1 2 2.39p
Rs 1 N3 0.34
L1 N3 2 30.423u
.ends 6033_7447785133_33u
*******
.subckt 6033_7447785147_47u 1 2
Rp 1 2 33526.9561318
Cp 1 2 2.43213501888p
Rs 1 N3 0.5
L1 N3 2 43.1174628648u
.ends 6033_7447785147_47u
*******
.subckt 6033_744778520_100u 1 2
Rp 1 2 61685.068896
Cp 1 2 2.81516160101p
Rs 1 N3 0.95
L1 N3 2 94.2316542955u
.ends 6033_744778520_100u
*******
.subckt 6050_7447786001_1u 1 2
Rp 1 2 2037.89824727
Cp 1 2 0.663634817p
Rs 1 N3 0.028
L1 N3 2 0.947508694023u
.ends 6050_7447786001_1u
*******
.subckt 6050_7447786002_2.2u 1 2
Rp 1 2 3873.12288939
Cp 1 2 0.888176917776p
Rs 1 N3 0.04
L1 N3 2 2.10110600258u
.ends 6050_7447786002_2.2u
*******
.subckt 6050_7447786004_4.7u 1 2
Rp 1 2 6482.96246684
Cp 1 2 2.13619859583p
Rs 1 N3 0.057
L1 N3 2 4.35584118762u
.ends 6050_7447786004_4.7u
*******
.subckt 6050_7447786006_6.8u 1 2
Rp 1 2 7197.76906562
Cp 1 2 2.28699835088p
Rs 1 N3 0.062
L1 N3 2 6.4423583094u
.ends 6050_7447786006_6.8u
*******
.subckt 6050_7447786008_8.2u 1 2
Rp 1 2 9510.40662457
Cp 1 2 2.2670543677p
Rs 1 N3 0.066
L1 N3 2 7.52568588616u
.ends 6050_7447786008_8.2u
*******
.subckt 6050_744778610_10u 1 2
Rp 1 2 10586.7671579
Cp 1 2 2.53999984512p
Rs 1 N3 0.074
L1 N3 2 8.34245072542u
.ends 6050_744778610_10u
*******
.subckt 6050_7447786122_22u 1 2
Rp 1 2 17374.7513097
Cp 1 2 5.64102666619p
Rs 1 N3 0.098
L1 N3 2 19.6300919502u
.ends 6050_7447786122_22u
*******
.subckt 6050_7447786147_47u 1 2
Rp 1 2 35068.1701337
Cp 1 2 5.79515468172p
Rs 1 N3 0.26
L1 N3 2 42.9111231439u
.ends 6050_7447786147_47u
*******
.subckt 7332_744778005_0.54u 1 2
Rp 1 2 1229.74139719
Cp 1 2 2.81710018376p
Rs 1 N3 0.0072
L1 N3 2 0.405637106674u
.ends 7332_744778005_0.54u
*******
.subckt 7332_7447789001_1u 1 2
Rp 1 2 2164.87869848
Cp 1 2 2.61396727902p
Rs 1 N3 0.01
L1 N3 2 0.772776226124u
.ends 7332_7447789001_1u
*******
.subckt 7332_744778001_1u 1 2
Rp 1 2 2166.12668275
Cp 1 2 2.47067045874p
Rs 1 N3 0.009
L1 N3 2 0.773397441523u
.ends 7332_744778001_1u
*******
.subckt 7332_7447783015_1.5u 1 2
Rp 1 2 1060
Cp 1 2 3.397p
Rs 1 N3 0.012
L1 N3 2 1.41u
.ends 7332_7447783015_1.5u
*******
.subckt 7332_7447789002_2.2u 1 2
Rp 1 2 5113.0951551
Cp 1 2 2.75488097451p
Rs 1 N3 0.019
L1 N3 2 2.0669826351u
.ends 7332_7447789002_2.2u
*******
.subckt 7332_744778002_2.2u 1 2
Rp 1 2 4984.65903378
Cp 1 2 2.66299907004p
Rs 1 N3 0.014
L1 N3 2 2.09435585344u
.ends 7332_744778002_2.2u
*******
.subckt 7332_7447783022_2.2u 1 2
Rp 1 2 1644
Cp 1 2 3.131p
Rs 1 N3 0.0155
L1 N3 2 2.11u
.ends 7332_7447783022_2.2u
*******
.subckt 7332_744778003_3.3u 1 2
Rp 1 2 6426.52613323
Cp 1 2 2.99661324441p
Rs 1 N3 0.024
L1 N3 2 2.56462716755u
.ends 7332_744778003_3.3u
*******
.subckt 7332_7447789003_3.3u 1 2
Rp 1 2 6967.01278729
Cp 1 2 2.34363124437p
Rs 1 N3 0.024
L1 N3 2 2.81530333037u
.ends 7332_7447789003_3.3u
*******
.subckt 7332_7447783033_3.3u 1 2
Rp 1 2 2339
Cp 1 2 3.477p
Rs 1 N3 0.018
L1 N3 2 2.88u
.ends 7332_7447783033_3.3u
*******
.subckt 7332_7447789004_4.7u 1 2
Rp 1 2 9174.29236527
Cp 1 2 3.00846976512p
Rs 1 N3 0.033
L1 N3 2 3.86514286773u
.ends 7332_7447789004_4.7u
*******
.subckt 7332_744778004_4.7u 1 2
Rp 1 2 8887.11646987
Cp 1 2 3.26091741837p
Rs 1 N3 0.042
L1 N3 2 4.06187686187u
.ends 7332_744778004_4.7u
*******
.subckt 7332_7447783047_4.7u 1 2
Rp 1 2 4208
Cp 1 2 3.56p
Rs 1 N3 0.027
L1 N3 2 4.08u
.ends 7332_7447783047_4.7u
*******
.subckt 7332_7447789006_6.8u 1 2
Rp 1 2 11163.6489624
Cp 1 2 3.1698604005p
Rs 1 N3 0.0415
L1 N3 2 5.82987393511u
.ends 7332_7447789006_6.8u
*******
.subckt 7332_7447783068_6.8u 1 2
Rp 1 2 5309
Cp 1 2 3.232p
Rs 1 N3 0.033
L1 N3 2 6.39u
.ends 7332_7447783068_6.8u
*******
.subckt 7332_74477810_10u 1 2
Rp 1 2 14371.7275969
Cp 1 2 3.06494111157p
Rs 1 N3 0.068
L1 N3 2 7.79780559887u
.ends 7332_74477810_10u
*******
.subckt 7332_744778910_10u 1 2
Rp 1 2 16852.2449006
Cp 1 2 2.7268024532p
Rs 1 N3 0.064
L1 N3 2 8.0668901277u
.ends 7332_744778910_10u
*******
.subckt 7332_7447783100_10u 1 2
Rp 1 2 8092
Cp 1 2 2.937p
Rs 1 N3 0.056
L1 N3 2 9.541u
.ends 7332_7447783100_10u
*******
.subckt 7332_744778112_12u 1 2
Rp 1 2 16520.2293361
Cp 1 2 3.43671378309p
Rs 1 N3 0.076
L1 N3 2 9.86176498616u
.ends 7332_744778112_12u
*******
.subckt 7332_7447789112_12u 1 2
Rp 1 2 19926.4041255
Cp 1 2 3.19462974993p
Rs 1 N3 0.076
L1 N3 2 10.341959258u
.ends 7332_7447789112_12u
*******
.subckt 7332_7447789115_15u 1 2
Rp 1 2 26979.0113761
Cp 1 2 2.95751468157p
Rs 1 N3 0.1
L1 N3 2 12.6691187155u
.ends 7332_7447789115_15u
*******
.subckt 7332_744778115_15u 1 2
Rp 1 2 22047.7802689
Cp 1 2 2.94868309515p
Rs 1 N3 0.1
L1 N3 2 13.1759854422u
.ends 7332_744778115_15u
*******
.subckt 7332_7447783150_15u 1 2
Rp 1 2 12813
Cp 1 2 3.463p
Rs 1 N3 0.068
L1 N3 2 13.88u
.ends 7332_7447783150_15u
*******
.subckt 7332_744778118_18u 1 2
Rp 1 2 23442.984673
Cp 1 2 3.33396069523p
Rs 1 N3 0.114
L1 N3 2 14.3694967628u
.ends 7332_744778118_18u
*******
.subckt 7332_7447789118_18u 1 2
Rp 1 2 32318.4705556
Cp 1 2 2.54642147041p
Rs 1 N3 0.114
L1 N3 2 16.2685632654u
.ends 7332_7447789118_18u
*******
.subckt 7332_744778122_22u 1 2
Rp 1 2 24860.2777908
Cp 1 2 3.71054637911p
Rs 1 N3 0.119
L1 N3 2 17.7891180195u
.ends 7332_744778122_22u
*******
.subckt 7332_7447783220_22u 1 2
Rp 1 2 18288
Cp 1 2 3.927p
Rs 1 N3 0.09
L1 N3 2 20.42u
.ends 7332_7447783220_22u
*******
.subckt 7332_7447789122_22u 1 2
Rp 1 2 33532.7850569
Cp 1 2 3.0576419453p
Rs 1 N3 0.119
L1 N3 2 20.6444606452u
.ends 7332_7447789122_22u
*******
.subckt 7332_7447789127_27u 1 2
Rp 1 2 37364.8490068
Cp 1 2 3.17982011113p
Rs 1 N3 0.13
L1 N3 2 23.0129196272u
.ends 7332_7447789127_27u
*******
.subckt 7332_744778127_27u 1 2
Rp 1 2 29087.5887631
Cp 1 2 3.4842205739p
Rs 1 N3 0.14
L1 N3 2 23.1463214499u
.ends 7332_744778127_27u
*******
.subckt 7332_744778133_33u 1 2
Rp 1 2 32451.612057
Cp 1 2 3.8300734141p
Rs 1 N3 0.153
L1 N3 2 25.3774240703u
.ends 7332_744778133_33u
*******
.subckt 7332_7447789133_33u 1 2
Rp 1 2 39404.9439766
Cp 1 2 3.54126090611p
Rs 1 N3 0.153
L1 N3 2 26.8716084055u
.ends 7332_7447789133_33u
*******
.subckt 7332_7447783330_33u 1 2
Rp 1 2 26459
Cp 1 2 4.227p
Rs 1 N3 0.138
L1 N3 2 30.89u
.ends 7332_7447783330_33u
*******
.subckt 7332_744778139_39u 1 2
Rp 1 2 41433.6642926
Cp 1 2 3.07597814933p
Rs 1 N3 0.214
L1 N3 2 31.098539109u
.ends 7332_744778139_39u
*******
.subckt 7332_7447789139_39u 1 2
Rp 1 2 34754.859201
Cp 1 2 3.46116451404p
Rs 1 N3 0.209
L1 N3 2 32.4605379645u
.ends 7332_7447789139_39u
*******
.subckt 7332_744778147_47u 1 2
Rp 1 2 48650.9889075
Cp 1 2 3.34473024276p
Rs 1 N3 0.315
L1 N3 2 39.1639576114u
.ends 7332_744778147_47u
*******
.subckt 7332_7447789147_47u 1 2
Rp 1 2 63191.9226458
Cp 1 2 3.41998431982p
Rs 1 N3 0.315
L1 N3 2 42.3770489237u
.ends 7332_7447789147_47u
*******
.subckt 7332_7447783470_47u 1 2
Rp 1 2 34357
Cp 1 2 4.3p
Rs 1 N3 0.18
L1 N3 2 43.58u
.ends 7332_7447783470_47u
*******
.subckt 7332_744778156_56u 1 2
Rp 1 2 54236.4427989
Cp 1 2 3.56528937344p
Rs 1 N3 0.322
L1 N3 2 46.7472808258u
.ends 7332_744778156_56u
*******
.subckt 7332_7447789156_56u 1 2
Rp 1 2 80877.7141423
Cp 1 2 3.08743856235p
Rs 1 N3 0.335
L1 N3 2 51.0054622523u
.ends 7332_7447789156_56u
*******
.subckt 7332_744778168_68u 1 2
Rp 1 2 59515.6102582
Cp 1 2 3.13894039646p
Rs 1 N3 0.417
L1 N3 2 57.6153789573u
.ends 7332_744778168_68u
*******
.subckt 7332_7447789168_68u 1 2
Rp 1 2 70531.1230274
Cp 1 2 3.20660212416p
Rs 1 N3 0.427
L1 N3 2 62.3263343297u
.ends 7332_7447789168_68u
*******
.subckt 7332_7447783680_68u 1 2
Rp 1 2 47333
Cp 1 2 4.393p
Rs 1 N3 0.26
L1 N3 2 65.94u
.ends 7332_7447783680_68u
*******
.subckt 7332_744778182_82u 1 2
Rp 1 2 73920.3213959
Cp 1 2 3.66660676379p
Rs 1 N3 0.479
L1 N3 2 72.7163371541u
.ends 7332_744778182_82u
*******
.subckt 7332_7447789182_82u 1 2
Rp 1 2 88537.3761503
Cp 1 2 3.47297926442p
Rs 1 N3 0.47
L1 N3 2 78.5446378433u
.ends 7332_7447789182_82u
*******
.subckt 7332_74477820_100u 1 2
Rp 1 2 65000
Cp 1 2 3.5p
Rs 1 N3 0.585
L1 N3 2 90u
.ends 7332_74477820_100u
*******
.subckt 7332_744778920_100u 1 2
Rp 1 2 101005.134156
Cp 1 2 3.44049203882p
Rs 1 N3 0.585
L1 N3 2 90.5473485736u
.ends 7332_744778920_100u
*******
.subckt 7332_744778212_120u 1 2
Rp 1 2 78183.3998498
Cp 1 2 3.10879750953p
Rs 1 N3 0.634
L1 N3 2 92.7530315334u
.ends 7332_744778212_120u
*******
.subckt 7332_7447783101_100u 1 2
Rp 1 2 59499
Cp 1 2 4.267p
Rs 1 N3 0.39
L1 N3 2 96.9u
.ends 7332_7447783101_100u
*******
.subckt 7332_7447789212_120u 1 2
Rp 1 2 120249.3167384
Cp 1 2 3.48227471573p
Rs 1 N3 0.563
L1 N3 2 104.788185426u
.ends 7332_7447789212_120u
*******
.subckt 7332_7447789215_150u 1 2
Rp 1 2 136237.960919
Cp 1 2 3.84852382952p
Rs 1 N3 0.72
L1 N3 2 127.718005681u
.ends 7332_7447789215_150u
*******
.subckt 7332_744778215_150u 1 2
Rp 1 2 90182.9907411
Cp 1 2 3.82610257368p
Rs 1 N3 0.72
L1 N3 2 128.618162736u
.ends 7332_744778215_150u
*******
.subckt 7332_7447783151_150u 1 2
Rp 1 2 80323
Cp 1 2 4.449p
Rs 1 N3 0.63
L1 N3 2 148.62u
.ends 7332_7447783151_150u
*******
.subckt 7332_744778218_180u 1 2
Rp 1 2 122686.047456
Cp 1 2 2.96881569994p
Rs 1 N3 0.96
L1 N3 2 153.788184817u
.ends 7332_744778218_180u
*******
.subckt 7332_7447789218_180u 1 2
Rp 1 2 121990.7268892
Cp 1 2 3.59620213037p
Rs 1 N3 0.96
L1 N3 2 155.387115339u
.ends 7332_7447789218_180u
*******
.subckt 7332_7447789222_220u 1 2
Rp 1 2 145290.519218
Cp 1 2 3.98898377328p
Rs 1 N3 1.35
L1 N3 2 178.2592594u
.ends 7332_7447789222_220u
*******
.subckt 7332_744778222_220u 1 2
Rp 1 2 144955.490273
Cp 1 2 3.83371324993p
Rs 1 N3 1.22
L1 N3 2 194.128533701u
.ends 7332_744778222_220u
*******
.subckt 7332_7447783221_220u 1 2
Rp 1 2 97034
Cp 1 2 4.72p
Rs 1 N3 0.87
L1 N3 2 216.71u
.ends 7332_7447783221_220u
*******
.subckt 7332_744778270_270u 1 2
Rp 1 2 147574.231316
Cp 1 2 4.4241022573p
Rs 1 N3 1.44
L1 N3 2 219.384019027u
.ends 7332_744778270_270u
*******
.subckt 7332_7447789270_270u 1 2
Rp 1 2 161634.517973
Cp 1 2 3.5539395336p
Rs 1 N3 1.47
L1 N3 2 249.40645638u
.ends 7332_7447789270_270u
*******
.subckt 7332_744778233_330u 1 2
Rp 1 2 190366.905413
Cp 1 2 3.82078679735p
Rs 1 N3 2.28
L1 N3 2 283.542394332u
.ends 7332_744778233_330u
*******
.subckt 7332_7447789233_330u 1 2
Rp 1 2 194710.510845
Cp 1 2 3.54039630514p
Rs 1 N3 2.28
L1 N3 2 301.724670852u
.ends 7332_7447789233_330u
*******
.subckt 7332_7447783331_330u 1 2
Rp 1 2 118446
Cp 1 2 5.0053p
Rs 1 N3 1.24
L1 N3 2 321.17u
.ends 7332_7447783331_330u
*******
.subckt 7332_744778239_390u 1 2
Rp 1 2 184242.489449
Cp 1 2 3.98514039572p
Rs 1 N3 2.49
L1 N3 2 324.897187206u
.ends 7332_744778239_390u
*******
.subckt 7332_7447789239_390u 1 2
Rp 1 2 207587.080246
Cp 1 2 3.66077620731p
Rs 1 N3 2.49
L1 N3 2 350.383943323u
.ends 7332_7447789239_390u
*******
.subckt 7332_74477824_470u 1 2
Rp 1 2 187991.752291
Cp 1 2 3.94647112544p
Rs 1 N3 2.6
L1 N3 2 402.122235065u
.ends 7332_74477824_470u
*******
.subckt 7332_744778924_470u 1 2
Rp 1 2 248636.618754
Cp 1 2 3.79414274243p
Rs 1 N3 2.6
L1 N3 2 408.480958848u
.ends 7332_744778924_470u
*******
.subckt 7332_74477830_1000u 1 2
Rp 1 2 124583.875664
Cp 1 2 9.625193217p
Rs 1 N3 5.57
L1 N3 2 418.147154636u
.ends 7332_74477830_1000u
*******
.subckt 7332_7447783471_470u 1 2
Rp 1 2 153394
Cp 1 2 5.1p
Rs 1 N3 1.78
L1 N3 2 457.06u
.ends 7332_7447783471_470u
*******
.subckt 7332_74477825_560u 1 2
Rp 1 2 184925.223731
Cp 1 2 4.11804015268p
Rs 1 N3 3
L1 N3 2 459.460469561u
.ends 7332_74477825_560u
*******
.subckt 7332_744778925_560u 1 2
Rp 1 2 301244.783132
Cp 1 2 3.35959221812p
Rs 1 N3 3
L1 N3 2 567.115841247u
.ends 7332_744778925_560u
*******
.subckt 7332_74477826_680u 1 2
Rp 1 2 210302.691304
Cp 1 2 4.02469121246p
Rs 1 N3 4.5
L1 N3 2 572.154405014u
.ends 7332_74477826_680u
*******
.subckt 7332_7447783681_680u 1 2
Rp 1 2 174162
Cp 1 2 5.219p
Rs 1 N3 2.52
L1 N3 2 641.24u
.ends 7332_7447783681_680u
*******
.subckt 7332_74477828_820u 1 2
Rp 1 2 372995.147279
Cp 1 2 4.41613646321p
Rs 1 N3 5.07
L1 N3 2 657.025953673u
.ends 7332_74477828_820u
*******
.subckt 7332_744778926_680u 1 2
Rp 1 2 373585.98853
Cp 1 2 3.83777523956p
Rs 1 N3 4.5
L1 N3 2 663.276647609u
.ends 7332_744778926_680u
*******
.subckt 7332_744778928_820u 1 2
Rp 1 2 597284.327437
Cp 1 2 3.69644017246p
Rs 1 N3 4.99
L1 N3 2 776.704667792u
.ends 7332_744778928_820u
*******
.subckt 7332_744778930_1000u 1 2
Rp 1 2 624396.631432
Cp 1 2 3.96080843446p
Rs 1 N3 5.57
L1 N3 2 908.1614785u
.ends 7332_744778930_1000u
*******
.subckt 7332_7447783102_1000u 1 2
Rp 1 2 226939
Cp 1 2 5.4977p
Rs 1 N3 4
L1 N3 2 950.14u
.ends 7332_7447783102_1000u
*******
.subckt 7345_7447773010_1u 1 2
Rp 1 2 552
Cp 1 2 3.126p
Rs 1 N3 0.0084
L1 N3 2 0.872u
.ends 7345_7447773010_1u
*******
.subckt 7345_744777001_1u 1 2
Rp 1 2 2428.067211
Cp 1 2 3.37078710741p
Rs 1 N3 0.0084
L1 N3 2 0.888631308826u
.ends 7345_744777001_1u
*******
.subckt 7345_7447779001_1u 1 2
Rp 1 2 2646.3028188
Cp 1 2 2.93181424014p
Rs 1 N3 0.01
L1 N3 2 0.953249649186u
.ends 7345_7447779001_1u
*******
.subckt 7345_74477790015_1.5u 1 2
Rp 1 2 3475.57841959
Cp 1 2 3.12984014451p
Rs 1 N3 0.015
L1 N3 2 1.49681672213u
.ends 7345_74477790015_1.5u
*******
.subckt 7345_744777002_2.2u 1 2
Rp 1 2 4447.62481375
Cp 1 2 3.0264444023p
Rs 1 N3 0.013
L1 N3 2 1.97916261562u
.ends 7345_744777002_2.2u
*******
.subckt 7345_7447773022_2.2u 1 2
Rp 1 2 1414
Cp 1 2 3.365p
Rs 1 N3 0.0125
L1 N3 2 2.008u
.ends 7345_7447773022_2.2u
*******
.subckt 7345_7447779002_2.2u 1 2
Rp 1 2 4374.75290382
Cp 1 2 3.53414711028p
Rs 1 N3 0.016
L1 N3 2 2.0226563278u
.ends 7345_7447779002_2.2u
*******
.subckt 7345_744777003_3.3u 1 2
Rp 1 2 5751.28754081
Cp 1 2 2.88912716099p
Rs 1 N3 0.025
L1 N3 2 2.53717040164u
.ends 7345_744777003_3.3u
*******
.subckt 7345_7447779003_3.3u 1 2
Rp 1 2 5748.82909593
Cp 1 2 2.68748396769p
Rs 1 N3 0.026
L1 N3 2 2.71820601429u
.ends 7345_7447779003_3.3u
*******
.subckt 7345_7447773033_3.3u 1 2
Rp 1 2 2136
Cp 1 2 3.187p
Rs 1 N3 0.0155
L1 N3 2 3.037u
.ends 7345_7447773033_3.3u
*******
.subckt 7345_744777004_4.7u 1 2
Rp 1 2 7181.46846934
Cp 1 2 4.74613294276p
Rs 1 N3 0.025
L1 N3 2 3.91390400368u
.ends 7345_744777004_4.7u
*******
.subckt 7345_7447779004_4.7u 1 2
Rp 1 2 7362.44264815
Cp 1 2 4.45138899616p
Rs 1 N3 0.028
L1 N3 2 4.03449474678u
.ends 7345_7447779004_4.7u
*******
.subckt 7345_7447773047_4.7u 1 2
Rp 1 2 3854
Cp 1 2 4.391p
Rs 1 N3 0.02
L1 N3 2 4.601u
.ends 7345_7447773047_4.7u
*******
.subckt 7345_7447779006_6.8u 1 2
Rp 1 2 9935.28889881
Cp 1 2 4.51363958015p
Rs 1 N3 0.033
L1 N3 2 5.50661603545u
.ends 7345_7447779006_6.8u
*******
.subckt 7345_7447773062_6.2u 1 2
Rp 1 2 5168
Cp 1 2 4.339p
Rs 1 N3 0.025
L1 N3 2 5.997u
.ends 7345_7447773062_6.2u
*******
.subckt 7345_7447779008_8.2u 1 2
Rp 1 2 12904.2197053
Cp 1 2 4.30943185861p
Rs 1 N3 0.047
L1 N3 2 7.74425370543u
.ends 7345_7447779008_8.2u
*******
.subckt 7345_74477710_10u 1 2
Rp 1 2 14381.9104507
Cp 1 2 4.71830999092p
Rs 1 N3 0.045
L1 N3 2 8.15133607688u
.ends 7345_74477710_10u
*******
.subckt 7345_744777910_10u 1 2
Rp 1 2 14923.8050022
Cp 1 2 4.35681550134p
Rs 1 N3 0.045
L1 N3 2 9.30399593124u
.ends 7345_744777910_10u
*******
.subckt 7345_7447773100_10u 1 2
Rp 1 2 9166
Cp 1 2 4.545p
Rs 1 N3 0.0375
L1 N3 2 10.406u
.ends 7345_7447773100_10u
*******
.subckt 7345_7447779112_12u 1 2
Rp 1 2 17359.8565677
Cp 1 2 4.70534602246p
Rs 1 N3 0.05
L1 N3 2 10.7587538076u
.ends 7345_7447779112_12u
*******
.subckt 7345_744777112_12u 1 2
Rp 1 2 16199.3519734
Cp 1 2 5.01854838019p
Rs 1 N3 0.054
L1 N3 2 10.8548790404u
.ends 7345_744777112_12u
*******
.subckt 7345_744777115_15u 1 2
Rp 1 2 20614.9376125
Cp 1 2 4.82966144472p
Rs 1 N3 0.07
L1 N3 2 13.2872063758u
.ends 7345_744777115_15u
*******
.subckt 7345_7447773150_15u 1 2
Rp 1 2 12187
Cp 1 2 4.461p
Rs 1 N3 0.053
L1 N3 2 13.36u
.ends 7345_7447773150_15u
*******
.subckt 7345_744777118_18u 1 2
Rp 1 2 19184.0823276
Cp 1 2 5.2698569186p
Rs 1 N3 0.08
L1 N3 2 14.0031324899u
.ends 7345_744777118_18u
*******
.subckt 7345_7447779115_15u 1 2
Rp 1 2 21289.9423556
Cp 1 2 4.64898874212p
Rs 1 N3 0.07
L1 N3 2 14.0553867045u
.ends 7345_7447779115_15u
*******
.subckt 7345_7447779118_18u 1 2
Rp 1 2 23352.4066309
Cp 1 2 4.83768050426p
Rs 1 N3 0.08
L1 N3 2 15.1365751407u
.ends 7345_7447779118_18u
*******
.subckt 7345_744777122_22u 1 2
Rp 1 2 25621.8097743
Cp 1 2 4.81862359532p
Rs 1 N3 0.09
L1 N3 2 17.312069208u
.ends 7345_744777122_22u
*******
.subckt 7345_7447779122_22u 1 2
Rp 1 2 26201.7154972
Cp 1 2 4.23269590731p
Rs 1 N3 0.09
L1 N3 2 19.6930183853u
.ends 7345_7447779122_22u
*******
.subckt 7345_7447773220_22u 1 2
Rp 1 2 18190
Cp 1 2 4.464p
Rs 1 N3 0.075
L1 N3 2 21.7u
.ends 7345_7447773220_22u
*******
.subckt 7345_744777127_27u 1 2
Rp 1 2 25969.5408515
Cp 1 2 6.30104455742p
Rs 1 N3 0.1172
L1 N3 2 21.9552246523u
.ends 7345_744777127_27u
*******
.subckt 7345_7447779127_27u 1 2
Rp 1 2 33172.6662422
Cp 1 2 5.73286736266p
Rs 1 N3 0.12
L1 N3 2 23.3493656033u
.ends 7345_7447779127_27u
*******
.subckt 7345_744777133_33u 1 2
Rp 1 2 31532.58464
Cp 1 2 5.54301558717p
Rs 1 N3 0.14
L1 N3 2 25.3587498061u
.ends 7345_744777133_33u
*******
.subckt 7345_7447779133_33u 1 2
Rp 1 2 33602.6479344
Cp 1 2 5.03887187495p
Rs 1 N3 0.14
L1 N3 2 27.5700648448u
.ends 7345_7447779133_33u
*******
.subckt 7345_7447773330_33u 1 2
Rp 1 2 23316
Cp 1 2 4.61p
Rs 1 N3 0.12
L1 N3 2 30.42u
.ends 7345_7447773330_33u
*******
.subckt 7345_744777139_39u 1 2
Rp 1 2 37085.9724851
Cp 1 2 6.12679559834p
Rs 1 N3 0.145
L1 N3 2 32.8697102392u
.ends 7345_744777139_39u
*******
.subckt 7345_7447779139_39u 1 2
Rp 1 2 42921.2869045
Cp 1 2 5.83277468758p
Rs 1 N3 0.145
L1 N3 2 34.4193355788u
.ends 7345_7447779139_39u
*******
.subckt 7345_744777147_47u 1 2
Rp 1 2 45128.6756745
Cp 1 2 5.51496715314p
Rs 1 N3 0.17
L1 N3 2 39.9201792108u
.ends 7345_744777147_47u
*******
.subckt 7345_7447779147_47u 1 2
Rp 1 2 27787
Cp 1 2 4.61p
Rs 1 N3 0.19
L1 N3 2 42.37u
.ends 7345_7447779147_47u
*******
.subckt 7345_7447773470_47u 1 2
Rp 1 2 35578
Cp 1 2 5.346p
Rs 1 N3 0.15
L1 N3 2 44.8u
.ends 7345_7447773470_47u
*******
.subckt 7345_744777156_56u 1 2
Rp 1 2 51644.788073
Cp 1 2 5.0594289911p
Rs 1 N3 0.207
L1 N3 2 45.13236412u
.ends 7345_744777156_56u
*******
.subckt 7345_7447779156_56u 1 2
Rp 1 2 58516.8805777
Cp 1 2 5.2026080755p
Rs 1 N3 0.228
L1 N3 2 47.5175594632u
.ends 7345_7447779156_56u
*******
.subckt 7345_744777168_68u 1 2
Rp 1 2 57243.6120012
Cp 1 2 5.25275598423p
Rs 1 N3 0.239
L1 N3 2 56.1067931323u
.ends 7345_744777168_68u
*******
.subckt 7345_7447773680_68u 1 2
Rp 1 2 40263
Cp 1 2 5.889p
Rs 1 N3 0.19
L1 N3 2 61.816u
.ends 7345_7447773680_68u
*******
.subckt 7345_7447779168_68u 1 2
Rp 1 2 68182.8335292
Cp 1 2 4.76346605562p
Rs 1 N3 0.239
L1 N3 2 63.6273713572u
.ends 7345_7447779168_68u
*******
.subckt 7345_744777182_82u 1 2
Rp 1 2 68149.3545963
Cp 1 2 5.0274195156p
Rs 1 N3 0.257
L1 N3 2 64.6145372775u
.ends 7345_744777182_82u
*******
.subckt 7345_7447779182_82u 1 2
Rp 1 2 84240.0560821
Cp 1 2 4.75892530446p
Rs 1 N3 0.25
L1 N3 2 78.6538851191u
.ends 7345_7447779182_82u
*******
.subckt 7345_74477720_100u 1 2
Rp 1 2 79138.4858104
Cp 1 2 5.30562429717p
Rs 1 N3 0.29
L1 N3 2 80.0836908931u
.ends 7345_74477720_100u
*******
.subckt 7345_744777920_100u 1 2
Rp 1 2 89819.0358469
Cp 1 2 5.08611447106p
Rs 1 N3 0.29
L1 N3 2 90.7869346393u
.ends 7345_744777920_100u
*******
.subckt 7345_7447773101_100u 1 2
Rp 1 2 48300
Cp 1 2 6.114p
Rs 1 N3 0.27
L1 N3 2 93.078u
.ends 7345_7447773101_100u
*******
.subckt 7345_744777212_120u 1 2
Rp 1 2 100252.361874
Cp 1 2 5.27084159388p
Rs 1 N3 0.4
L1 N3 2 100.825421147u
.ends 7345_744777212_120u
*******
.subckt 7345_7447779212_120u 1 2
Rp 1 2 99257.6176478
Cp 1 2 5.24579465954p
Rs 1 N3 0.396
L1 N3 2 101.430158271u
.ends 7345_7447779212_120u
*******
.subckt 7345_744777215_150u 1 2
Rp 1 2 127685.790337
Cp 1 2 6.22006520702p
Rs 1 N3 0.66
L1 N3 2 122.858072284u
.ends 7345_744777215_150u
*******
.subckt 7345_7447779215_150u 1 2
Rp 1 2 126805.687293
Cp 1 2 5.35261473p
Rs 1 N3 0.529
L1 N3 2 137.055444894u
.ends 7345_7447779215_150u
*******
.subckt 7345_7447773151_150u 1 2
Rp 1 2 70802
Cp 1 2 6.463p
Rs 1 N3 0.41
L1 N3 2 144.5u
.ends 7345_7447773151_150u
*******
.subckt 7345_744777218_180u 1 2
Rp 1 2 114582.946626
Cp 1 2 5.53393291606p
Rs 1 N3 0.68
L1 N3 2 151.807099498u
.ends 7345_744777218_180u
*******
.subckt 7345_7447779218_180u 1 2
Rp 1 2 169631.359763
Cp 1 2 5.14698329059p
Rs 1 N3 0.603
L1 N3 2 162.221220598u
.ends 7345_7447779218_180u
*******
.subckt 7345_744777222_220u 1 2
Rp 1 2 162801.89931
Cp 1 2 5.43777181379p
Rs 1 N3 0.92
L1 N3 2 181.49166338u
.ends 7345_744777222_220u
*******
.subckt 7345_7447779222_220u 1 2
Rp 1 2 178284.450317
Cp 1 2 5.33528144763p
Rs 1 N3 0.92
L1 N3 2 185.690752965u
.ends 7345_7447779222_220u
*******
.subckt 7345_7447773221_220u 1 2
Rp 1 2 76374
Cp 1 2 6.216p
Rs 1 N3 0.64
L1 N3 2 213u
.ends 7345_7447773221_220u
*******
.subckt 7345_744777270_270u 1 2
Rp 1 2 196257.14623
Cp 1 2 5.60320567816p
Rs 1 N3 0.97
L1 N3 2 237.051562825u
.ends 7345_744777270_270u
*******
.subckt 7345_7447779270_270u 1 2
Rp 1 2 183606.401985
Cp 1 2 5.58950089371p
Rs 1 N3 1.09
L1 N3 2 240.787230442u
.ends 7345_7447779270_270u
*******
.subckt 7345_744777233_330u 1 2
Rp 1 2 118697.299222
Cp 1 2 5.63076805756p
Rs 1 N3 1.15
L1 N3 2 255.586412817u
.ends 7345_744777233_330u
*******
.subckt 7345_7447779233_330u 1 2
Rp 1 2 157498.120922
Cp 1 2 5.28214190974p
Rs 1 N3 1.15
L1 N3 2 284.452816324u
.ends 7345_7447779233_330u
*******
.subckt 7345_7447773331_330u 1 2
Rp 1 2 116602
Cp 1 2 6.216p
Rs 1 N3 0.9
L1 N3 2 318u
.ends 7345_7447773331_330u
*******
.subckt 7345_744777239_390u 1 2
Rp 1 2 181977.786297
Cp 1 2 5.39201947666p
Rs 1 N3 1.25
L1 N3 2 330.180475498u
.ends 7345_744777239_390u
*******
.subckt 7345_7447779239_390u 1 2
Rp 1 2 210937.586684
Cp 1 2 5.22562974371p
Rs 1 N3 1.4
L1 N3 2 345.286258765u
.ends 7345_7447779239_390u
*******
.subckt 7345_74477724_470u 1 2
Rp 1 2 211485.011889
Cp 1 2 5.89682390032p
Rs 1 N3 1.6
L1 N3 2 406.405191616u
.ends 7345_74477724_470u
*******
.subckt 7345_744777924_470u 1 2
Rp 1 2 244548.076127
Cp 1 2 6.54965252578p
Rs 1 N3 1.6
L1 N3 2 436.730523269u
.ends 7345_744777924_470u
*******
.subckt 7345_74477725_560u 1 2
Rp 1 2 221658.160265
Cp 1 2 6.1688290058p
Rs 1 N3 1.72
L1 N3 2 460.193784526u
.ends 7345_74477725_560u
*******
.subckt 7345_7447773471_470u 1 2
Rp 1 2 137529
Cp 1 2 6.974p
Rs 1 N3 1.36
L1 N3 2 468u
.ends 7345_7447773471_470u
*******
.subckt 7345_744777925_560u 1 2
Rp 1 2 262369.520347
Cp 1 2 5.59197086429p
Rs 1 N3 1.72
L1 N3 2 483.734943366u
.ends 7345_744777925_560u
*******
.subckt 7345_74477726_680u 1 2
Rp 1 2 230392.597719
Cp 1 2 6.20727965463p
Rs 1 N3 2.6
L1 N3 2 565.122792057u
.ends 7345_74477726_680u
*******
.subckt 7345_744777926_680u 1 2
Rp 1 2 273721.142891
Cp 1 2 5.63004137531p
Rs 1 N3 2.6
L1 N3 2 582.603956244u
.ends 7345_744777926_680u
*******
.subckt 7345_7447773681_680u 1 2
Rp 1 2 147765
Cp 1 2 7.154p
Rs 1 N3 1.95
L1 N3 2 656u
.ends 7345_7447773681_680u
*******
.subckt 7345_74477728_820u 1 2
Rp 1 2 324901.854346
Cp 1 2 6.41419541325p
Rs 1 N3 3
L1 N3 2 668.728777469u
.ends 7345_74477728_820u
*******
.subckt 7345_744777928_820u 1 2
Rp 1 2 307854.062137
Cp 1 2 6.06252057637p
Rs 1 N3 2.96
L1 N3 2 726.765626894u
.ends 7345_744777928_820u
*******
.subckt 7345_74477730_1000u 1 2
Rp 1 2 385124.331896
Cp 1 2 5.86126999151p
Rs 1 N3 3.27
L1 N3 2 788.749706864u
.ends 7345_74477730_1000u
*******
.subckt 7345_744777930_1000u 1 2
Rp 1 2 443864.014531
Cp 1 2 5.53950555762p
Rs 1 N3 3.27
L1 N3 2 894.357609262u
.ends 7345_744777930_1000u
*******
.subckt 7345_7447773102_1000u 1 2
Rp 1 2 260130
Cp 1 2 7.276p
Rs 1 N3 2.85
L1 N3 2 976u
.ends 7345_7447773102_1000u
*******
