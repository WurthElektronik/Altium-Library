**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Shielded Coupled Inductor
* Matchcode:              WE-TDC 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 8018_744894300033_0.33u  1  2  3  4  PARAMS:
+  Cww=0.485p
+  Rp1=763
+  Cp1=1.62p
+  Lp1=0.21u
+  Rp2=763
+  Cp2=1.62p
+  Lp2=0.21u
+  RDC1=0.0111
+  RDC2=0.0111
+  K=0.813
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_744894300068_0.68u  1  2  3  4  PARAMS:
+  Cww=1.2175p
+  Rp1=1283.06
+  Cp1=1.52p
+  Lp1=0.45u
+  Rp2=1283.06
+  Cp2=1.52p
+  Lp2=0.45u
+  RDC1=0.0163
+  RDC2=0.0163
+  K=0.904
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430010_1u  1  2  3  4  PARAMS:
+  Cww=1.6225p
+  Rp1=1948.86
+  Cp1=1.81p
+  Lp1=0.7u
+  Rp2=1948.86
+  Cp2=1.81p
+  Lp2=0.7u
+  RDC1=0.0222
+  RDC2=0.0222
+  K=0.93
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430022_2.2u  1  2  3  4  PARAMS:
+  Cww=2.1975p
+  Rp1=3806.4
+  Cp1=1.89p
+  Lp1=1.53u
+  Rp2=3806.4
+  Cp2=1.89p
+  Lp2=1.53u
+  RDC1=0.0495
+  RDC2=0.0495
+  K=0.477
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430027_2.7u  1  2  3  4  PARAMS:
+  Cww=3.4525p
+  Rp1=4838.14
+  Cp1=2.29p
+  Lp1=1.98u
+  Rp2=4838.14
+  Cp2=2.29p
+  Lp2=1.98u
+  RDC1=0.0695
+  RDC2=0.0695
+  K=0.962
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430039_3.9u  1  2  3  4  PARAMS:
+  Cww=3.905p
+  Rp1=5329.33
+  Cp1=2.36p
+  Lp1=2.66u
+  Rp2=5329.33
+  Cp2=2.36p
+  Lp2=2.66u
+  RDC1=0.082
+  RDC2=0.082
+  K=0.976
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430056_5.6u  1  2  3  4  PARAMS:
+  Cww=5.7725p
+  Rp1=7670.19
+  Cp1=2.2p
+  Lp1=4.34u
+  Rp2=7670.19
+  Cp2=2.2p
+  Lp2=4.34u
+  RDC1=0.114
+  RDC2=0.114
+  K=0.997
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430100_10u  1  2  3  4  PARAMS:
+  Cww=5.8025p
+  Rp1=11623.01
+  Cp1=2.17p
+  Lp1=7.32u
+  Rp2=11623.01
+  Cp2=2.17p
+  Lp2=7.32u
+  RDC1=0.19
+  RDC2=0.19
+  K=0.984
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430120_12u  1  2  3  4  PARAMS:
+  Cww=6.195p
+  Rp1=11.97
+  Cp1=2.49p
+  Lp1=8.4u
+  Rp2=11.97
+  Cp2=2.49p
+  Lp2=8.4u
+  RDC1=0.202
+  RDC2=0.202
+  K=0.985
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430150_15u  1  2  3  4  PARAMS:
+  Cww=6.1975p
+  Rp1=15148.49
+  Cp1=2.15p
+  Lp1=11.26u
+  Rp2=15148.49
+  Cp2=2.15p
+  Lp2=11.26u
+  RDC1=0.262
+  RDC2=0.262
+  K=0.981
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8018_74489430180_18u  1  2  3  4  PARAMS:
+  Cww=7.5125p
+  Rp1=15346.68
+  Cp1=2.43p
+  Lp1=13.42u
+  Rp2=15346.68
+  Cp2=2.43p
+  Lp2=13.42u
+  RDC1=0.345
+  RDC2=0.345
+  K=0.987
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_744894400039_0.39u  1  2  3  4  PARAMS:
+  Cww=0.2625p
+  Rp1=924.87
+  Cp1=1.12p
+  Lp1=0.26u
+  Rp2=924.87
+  Cp2=1.12p
+  Lp2=0.26u
+  RDC1=0.0116
+  RDC2=0.0116
+  K=0.84
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_744894400082_0.82u  1  2  3  4  PARAMS:
+  Cww=1.115p
+  Rp1=1715.37
+  Cp1=1.36p
+  Lp1=0.57u
+  Rp2=1715.37
+  Cp2=1.36p
+  Lp2=0.57u
+  RDC1=0.0159
+  RDC2=0.0159
+  K=0.93
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440012_1.2u  1  2  3  4  PARAMS:
+  Cww=1.995p
+  Rp1=2576.03
+  Cp1=1.62p
+  Lp1=1.05u
+  Rp2=2576.03
+  Cp2=1.62p
+  Lp2=1.05u
+  RDC1=0.0202
+  RDC2=0.0202
+  K=0.954
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440018_1.8u  1  2  3  4  PARAMS:
+  Cww=1.8625p
+  Rp1=3094.71
+  Cp1=1.71p
+  Lp1=1.68u
+  Rp2=3094.71
+  Cp2=1.71p
+  Lp2=1.68u
+  RDC1=0.0255
+  RDC2=0.0255
+  K=0.979
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440027_2.7u  1  2  3  4  PARAMS:
+  Cww=3.9225p
+  Rp1=4176.26
+  Cp1=3.13p
+  Lp1=2.05u
+  Rp2=4176.26
+  Cp2=3.13p
+  Lp2=2.05u
+  RDC1=0.0345
+  RDC2=0.0345
+  K=0.954
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440036_3.6u  1  2  3  4  PARAMS:
+  Cww=3.4775p
+  Rp1=5788.12
+  Cp1=3.41p
+  Lp1=2.95u
+  Rp2=5788.12
+  Cp2=3.41p
+  Lp2=2.95u
+  RDC1=0.047
+  RDC2=0.047
+  K=0.941
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440047_4.7u  1  2  3  4  PARAMS:
+  Cww=4.7775p
+  Rp1=5491.59
+  Cp1=3.91p
+  Lp1=2.95u
+  Rp2=5491.59
+  Cp2=3.91p
+  Lp2=2.95u
+  RDC1=0.0545
+  RDC2=0.0545
+  K=0.973
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440120_12u  1  2  3  4  PARAMS:
+  Cww=10.53p
+  Rp1=10897.48
+  Cp1=5.06p
+  Lp1=9.7u
+  Rp2=10897.48
+  Cp2=5.06p
+  Lp2=9.7u
+  RDC1=0.117
+  RDC2=0.117
+  K=0.652
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440150_15u  1  2  3  4  PARAMS:
+  Cww=6.245p
+  Rp1=11343.48
+  Cp1=5.23p
+  Lp1=12.14u
+  Rp2=11343.48
+  Cp2=5.23p
+  Lp2=12.14u
+  RDC1=0.165
+  RDC2=0.165
+  K=0.981
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440180_18u  1  2  3  4  PARAMS:
+  Cww=8.58p
+  Rp1=15599.47
+  Cp1=5.29p
+  Lp1=15.73u
+  Rp2=15599.47
+  Cp2=5.29p
+  Lp2=15.73u
+  RDC1=0.179
+  RDC2=0.179
+  K=0.972
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
.subckt 8038_74489440220_22u  1  2  3  4  PARAMS:
+  Cww=12.9825p
+  Rp1=17240.33
+  Cp1=4.81p
+  Lp1=18.11u
+  Rp2=17240.33
+  Cp2=4.81p
+  Lp2=18.11u
+  RDC1=0.203
+  RDC2=0.203
+  K=0.988
C_C1  2  1    {Cww/2}
R_R50  2  1  5000g
C_C2  3  4    {Cww/2}
C_C5  3  2    {Cp1}
R_R1  3  N05454    {RDC1}
R_R2  3  2    {Rp1}
L_L1  N05454  2    {Lp1}
L_L2  N05750  1    {Lp2}
C_C6  4  1    {Cp2}
R_R3  4  1    {Rp2}
R_R4  4  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******
