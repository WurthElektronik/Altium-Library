**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  SMT Power Inductor
* Matchcode:              WE-LQS
* Library Type:           LTspice
* Version:                rev23a
* Created/modified by:    Ella
* Date and Time:          7/24/2023
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2023 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************
.subckt 2010_74404020010_1u 1 2
Rp 1 2 1870
Cp 1 2 1.129p
Rs 1 N3 0.094
L1 N3 2 0.724u
.ends 2010_74404020010_1u
*******
.subckt 2010_74404020015_1.5u 1 2
Rp 1 2 3137
Cp 1 2 1.093p
Rs 1 N3 0.147
L1 N3 2 1.24u
.ends 2010_74404020015_1.5u
*******
.subckt 2010_74404020022_2.2u 1 2
Rp 1 2 4597
Cp 1 2 1.191p
Rs 1 N3 0.225
L1 N3 2 1.789u
.ends 2010_74404020022_2.2u
*******
.subckt 2010_74404020033_3.3u 1 2
Rp 1 2 5074
Cp 1 2 1.396p
Rs 1 N3 0.275
L1 N3 2 3.148u
.ends 2010_74404020033_3.3u
*******
.subckt 2010_74404020047_4.7u 1 2
Rp 1 2 6490
Cp 1 2 1.338p
Rs 1 N3 0.41
L1 N3 2 4.013u
.ends 2010_74404020047_4.7u
*******
.subckt 2010_74404020068_6.8u 1 2
Rp 1 2 9099
Cp 1 2 1.346p
Rs 1 N3 0.7
L1 N3 2 6.754u
.ends 2010_74404020068_6.8u
*******
.subckt 2010_74404020100_10u 1 2
Rp 1 2 10056
Cp 1 2 1.922p
Rs 1 N3 0.86
L1 N3 2 9.062u
.ends 2010_74404020100_10u
*******
.subckt 2010_744040200016_0.16u 1 2
Rp 1 2 425
Cp 1 2 0.67p
Rs 1 N3 0.025
L1 N3 2 0.13u
.ends 2010_744040200016_0.16u
*******
.subckt 2010_744040200033_0.33u 1 2
Rp 1 2 735
Cp 1 2 0.747p
Rs 1 N3 0.034
L1 N3 2 0.288u
.ends 2010_744040200033_0.33u
*******
.subckt 2010_744040200047_0.47u 1 2
Rp 1 2 1157
Cp 1 2 0.86p
Rs 1 N3 0.047
L1 N3 2 0.365u
.ends 2010_744040200047_0.47u
*******
.subckt 2010_744040200068_0.68u 1 2
Rp 1 2 1521
Cp 1 2 1.254p
Rs 1 N3 0.064
L1 N3 2 0.501u
.ends 2010_744040200068_0.68u
*******
.subckt 2512_74404024010_1u 1 2
Rp 1 2 1700
Cp 1 2 1.34p
Rs 1 N3 0.036
L1 N3 2 0.789u
.ends 2512_74404024010_1u
*******
.subckt 2512_74404024015_1.5u 1 2
Rp 1 2 3236
Cp 1 2 0.869p
Rs 1 N3 0.065
L1 N3 2 1.302u
.ends 2512_74404024015_1.5u
*******
.subckt 2512_74404024022_2.2u 1 2
Rp 1 2 3570
Cp 1 2 2.07p
Rs 1 N3 0.08
L1 N3 2 1.7u
.ends 2512_74404024022_2.2u
*******
.subckt 2512_74404024033_3.3u 1 2
Rp 1 2 4630
Cp 1 2 2.25p
Rs 1 N3 0.12
L1 N3 2 2.9u
.ends 2512_74404024033_3.3u
*******
.subckt 2512_74404024047_4.7u 1 2
Rp 1 2 5220
Cp 1 2 1.56p
Rs 1 N3 0.173
L1 N3 2 4.57u
.ends 2512_74404024047_4.7u
*******
.subckt 2512_74404024068_6.8u 1 2
Rp 1 2 8630
Cp 1 2 2.4p
Rs 1 N3 0.3
L1 N3 2 6.59u
.ends 2512_74404024068_6.8u
*******
.subckt 2512_74404024100_10u 1 2
Rp 1 2 11070
Cp 1 2 2.14p
Rs 1 N3 0.43
L1 N3 2 8.87u
.ends 2512_74404024100_10u
*******
.subckt 2512_74404024150_15u 1 2
Rp 1 2 15522
Cp 1 2 1.5p
Rs 1 N3 0.82
L1 N3 2 17.13u
.ends 2512_74404024150_15u
*******
.subckt 2512_74404024180_18u 1 2
Rp 1 2 19400
Cp 1 2 2.33p
Rs 1 N3 0.83
L1 N3 2 15.7u
.ends 2512_74404024180_18u
*******
.subckt 2512_74404024220_22u 1 2
Rp 1 2 19400
Cp 1 2 2.4p
Rs 1 N3 0.91
L1 N3 2 21.6u
.ends 2512_74404024220_22u
*******
.subckt 2512_74404024330_33u 1 2
Rp 1 2 22500
Cp 1 2 1.45p
Rs 1 N3 1.53
L1 N3 2 40.5u
.ends 2512_74404024330_33u
*******
.subckt 2512_74404024470_47u 1 2
Rp 1 2 27000
Cp 1 2 1.66p
Rs 1 N3 1.65
L1 N3 2 56.3u
.ends 2512_74404024470_47u
*******
.subckt 2512_74404024680_68u 1 2
Rp 1 2 40100
Cp 1 2 2.23p
Rs 1 N3 2.4
L1 N3 2 78.5u
.ends 2512_74404024680_68u
*******
.subckt 2512_744040240016_0.16u 1 2
Rp 1 2 551.71
Cp 1 2 0.274p
Rs 1 N3 0.016
L1 N3 2 0.149u
.ends 2512_744040240016_0.16u
*******
.subckt 2512_744040240047_0.47u 1 2
Rp 1 2 1500
Cp 1 2 0.967p
Rs 1 N3 0.032
L1 N3 2 0.387u
.ends 2512_744040240047_0.47u
*******
.subckt 2512_744040240068_0.68u 1 2
Rp 1 2 1880
Cp 1 2 1.41p
Rs 1 N3 0.035
L1 N3 2 0.528u
.ends 2512_744040240068_0.68u
*******
.subckt 3015_74404032010_1u 1 2
Rp 1 2 1774.55518
Cp 1 2 1.7197657p
Rs 1 N3 0.033
L1 N3 2 0.849730568u
.ends 3015_74404032010_1u
*******
.subckt 3015_74404032015_1.5u 1 2
Rp 1 2 2250
Cp 1 2 1.97604444p
Rs 1 N3 0.04
L1 N3 2 1.2613888u
.ends 3015_74404032015_1.5u
*******
.subckt 3015_74404032022_2.2u 1 2
Rp 1 2 2946
Cp 1 2 1.203p
Rs 1 N3 0.05
L1 N3 2 1.751u
.ends 3015_74404032022_2.2u
*******
.subckt 3015_74404032033_3.3u 1 2
Rp 1 2 4117
Cp 1 2 1.80801396p
Rs 1 N3 0.07
L1 N3 2 2.54753468u
.ends 3015_74404032033_3.3u
*******
.subckt 3015_74404032047_4.7u 1 2
Rp 1 2 5434
Cp 1 2 2.19p
Rs 1 N3 0.096
L1 N3 2 4.173u
.ends 3015_74404032047_4.7u
*******
.subckt 3015_74404032068_6.8u 1 2
Rp 1 2 6025
Cp 1 2 1.3p
Rs 1 N3 0.12
L1 N3 2 6.784u
.ends 3015_74404032068_6.8u
*******
.subckt 3015_74404032100_10u 1 2
Rp 1 2 8884
Cp 1 2 3.2p
Rs 1 N3 0.23
L1 N3 2 8.05u
.ends 3015_74404032100_10u
*******
.subckt 3015_74404032101_100u 1 2
Rp 1 2 43750
Cp 1 2 2.5p
Rs 1 N3 1.9
L1 N3 2 115u
.ends 3015_74404032101_100u
*******
.subckt 3015_74404032150_15u 1 2
Rp 1 2 10800
Cp 1 2 3.46p
Rs 1 N3 0.3
L1 N3 2 12.97u
.ends 3015_74404032150_15u
*******
.subckt 3015_74404032220_22u 1 2
Rp 1 2 17435
Cp 1 2 1.4p
Rs 1 N3 0.45
L1 N3 2 20.8u
.ends 3015_74404032220_22u
*******
.subckt 3015_74404032330_33u 1 2
Rp 1 2 25400
Cp 1 2 2.1p
Rs 1 N3 0.911
L1 N3 2 28.9u
.ends 3015_74404032330_33u
*******
.subckt 3015_74404032470_47u 1 2
Rp 1 2 28731
Cp 1 2 2.9p
Rs 1 N3 1.05
L1 N3 2 41.8u
.ends 3015_74404032470_47u
*******
.subckt 3015_74404032680_68u 1 2
Rp 1 2 30860
Cp 1 2 2.06p
Rs 1 N3 1.6
L1 N3 2 76u
.ends 3015_74404032680_68u
*******
.subckt 3015_744040320047_0.47u 1 2
Rp 1 2 893.048
Cp 1 2 0.609p
Rs 1 N3 0.018
L1 N3 2 0.4061u
.ends 3015_744040320047_0.47u
*******
.subckt 4012_74404041010_1u 1 2
Rp 1 2 1846
Cp 1 2 0.939618p
Rs 1 N3 0.041
L1 N3 2 0.978u
.ends 4012_74404041010_1u
*******
.subckt 4012_74404041033_3.3u 1 2
Rp 1 2 3665
Cp 1 2 1.786p
Rs 1 N3 0.069
L1 N3 2 3.04u
.ends 4012_74404041033_3.3u
*******
.subckt 4012_74404041047_4.7u 1 2
Rp 1 2 4302
Cp 1 2 1.228p
Rs 1 N3 0.091
L1 N3 2 4.614u
.ends 4012_74404041047_4.7u
*******
.subckt 4012_74404041100_10u 1 2
Rp 1 2 7690
Cp 1 2 1.352p
Rs 1 N3 0.168
L1 N3 2 9.355u
.ends 4012_74404041100_10u
*******
.subckt 4012_74404041101_100u 1 2
Rp 1 2 30010
Cp 1 2 2.67p
Rs 1 N3 1.697
L1 N3 2 79.659u
.ends 4012_74404041101_100u
*******
.subckt 4012_74404041220_22u 1 2
Rp 1 2 13535
Cp 1 2 2.206p
Rs 1 N3 0.38
L1 N3 2 20.804u
.ends 4012_74404041220_22u
*******
.subckt 4012_74404041330_33u 1 2
Rp 1 2 16475
Cp 1 2 3.245p
Rs 1 N3 0.628
L1 N3 2 33.799u
.ends 4012_74404041330_33u
*******
.subckt 4012_74404041470_47u 1 2
Rp 1 2 23546
Cp 1 2 1.626p
Rs 1 N3 0.987
L1 N3 2 40.606u
.ends 4012_74404041470_47u
*******
.subckt 4012_74404041680_68u 1 2
Rp 1 2 28590
Cp 1 2 3.298p
Rs 1 N3 1.495
L1 N3 2 64.172u
.ends 4012_74404041680_68u
*******
.subckt 4012_744040410047_0.47u 1 2
Rp 1 2 689.207
Cp 1 2 0.480332p
Rs 1 N3 0.028
L1 N3 2 0.39093u
.ends 4012_744040410047_0.47u
*******
.subckt 4018_74404042010_1u 1 2
Rp 1 2 2364
Cp 1 2 1.213p
Rs 1 N3 0.027
L1 N3 2 0.999u
.ends 4018_74404042010_1u
*******
.subckt 4018_74404042015_1.5u 1 2
Rp 1 2 2627.9691
Cp 1 2 2.4928823p
Rs 1 N3 0.031
L1 N3 2 1.1246677u
.ends 4018_74404042015_1.5u
*******
.subckt 4018_74404042022_2.2u 1 2
Rp 1 2 3751.81556
Cp 1 2 2.5502999p
Rs 1 N3 0.042
L1 N3 2 1.8152807u
.ends 4018_74404042022_2.2u
*******
.subckt 4018_74404042033_3.3u 1 2
Rp 1 2 4325
Cp 1 2 2.257p
Rs 1 N3 0.055
L1 N3 2 3.172u
.ends 4018_74404042033_3.3u
*******
.subckt 4018_74404042047_4.7u 1 2
Rp 1 2 4582.6134
Cp 1 2 3.17959888p
Rs 1 N3 0.07
L1 N3 2 2.56204594u
.ends 4018_74404042047_4.7u
*******
.subckt 4018_74404042068_6.8u 1 2
Rp 1 2 6810.11761666667
Cp 1 2 2.93005643333333p
Rs 1 N3 0.098
L1 N3 2 5.4764569u
.ends 4018_74404042068_6.8u
*******
.subckt 4018_74404042100_10u 1 2
Rp 1 2 8513
Cp 1 2 2.268p
Rs 1 N3 0.15
L1 N3 2 9.042u
.ends 4018_74404042100_10u
*******
.subckt 4018_74404042101_100u 1 2
Rp 1 2 37616
Cp 1 2 2.947p
Rs 1 N3 1.43
L1 N3 2 91.193u
.ends 4018_74404042101_100u
*******
.subckt 4018_74404042150_15u 1 2
Rp 1 2 12553.3354
Cp 1 2 3.7005652p
Rs 1 N3 0.21
L1 N3 2 13.2308762u
.ends 4018_74404042150_15u
*******
.subckt 4018_74404042151_150u 1 2
Rp 1 2 60644
Cp 1 2 2.389p
Rs 1 N3 2.853
L1 N3 2 142.134u
.ends 4018_74404042151_150u
*******
.subckt 4018_74404042220_22u 1 2
Rp 1 2 15110.7838
Cp 1 2 4.36802208p
Rs 1 N3 0.29
L1 N3 2 18.2547578u
.ends 4018_74404042220_22u
*******
.subckt 4018_74404042221_220u 1 2
Rp 1 2 80520.6622
Cp 1 2 4.33334338p
Rs 1 N3 3.45
L1 N3 2 187.628388u
.ends 4018_74404042221_220u
*******
.subckt 4018_74404042330_33u 1 2
Rp 1 2 21390
Cp 1 2 2.554p
Rs 1 N3 0.46
L1 N3 2 29.071u
.ends 4018_74404042330_33u
*******
.subckt 4018_74404042331_330u 1 2
Rp 1 2 106007
Cp 1 2 3.584p
Rs 1 N3 5.3
L1 N3 2 305.113u
.ends 4018_74404042331_330u
*******
.subckt 4018_74404042470_47u 1 2
Rp 1 2 24493.3326
Cp 1 2 4.50042068p
Rs 1 N3 0.62
L1 N3 2 41.8222436u
.ends 4018_74404042470_47u
*******
.subckt 4018_74404042680_68u 1 2
Rp 1 2 29329.2486
Cp 1 2 5.61248904p
Rs 1 N3 0.84
L1 N3 2 61.3959988u
.ends 4018_74404042680_68u
*******
.subckt 4018_744040420033_0.33u 1 2
Rp 1 2 688
Cp 1 2 0.538976p
Rs 1 N3 0.013
L1 N3 2 0.283185u
.ends 4018_744040420033_0.33u
*******
.subckt 4025_74404043010A_1u 1 2
Rp 1 2 1430
Cp 1 2 1.37p
Rs 1 N3 0.014
L1 N3 2 0.695u
.ends 4025_74404043010A_1u
*******
.subckt 4025_74404043022A_2.2u 1 2
Rp 1 2 3300
Cp 1 2 1.535p
Rs 1 N3 0.023
L1 N3 2 1.464u
.ends 4025_74404043022A_2.2u
*******
.subckt 4025_74404043033A_3.3u 1 2
Rp 1 2 4750
Cp 1 2 1.78p
Rs 1 N3 0.033
L1 N3 2 2.48u
.ends 4025_74404043033A_3.3u
*******
.subckt 4025_74404043047A_4.7u 1 2
Rp 1 2 6060
Cp 1 2 1.835p
Rs 1 N3 0.046
L1 N3 2 3.67u
.ends 4025_74404043047A_4.7u
*******
.subckt 4025_74404043100A_10u 1 2
Rp 1 2 12650
Cp 1 2 1.92p
Rs 1 N3 0.089
L1 N3 2 7.73u
.ends 4025_74404043100A_10u
*******
.subckt 4025_74404043101A_100u 1 2
Rp 1 2 88400
Cp 1 2 2.43p
Rs 1 N3 1.043
L1 N3 2 87.7u
.ends 4025_74404043101A_100u
*******
.subckt 4025_74404043150A_15u 1 2
Rp 1 2 15700
Cp 1 2 2.3p
Rs 1 N3 0.132
L1 N3 2 11.78u
.ends 4025_74404043150A_15u
*******
.subckt 4025_74404043151A_150u 1 2
Rp 1 2 135800
Cp 1 2 2.36p
Rs 1 N3 1.634
L1 N3 2 125.3u
.ends 4025_74404043151A_150u
*******
.subckt 4025_74404043220A_22u 1 2
Rp 1 2 26600
Cp 1 2 2p
Rs 1 N3 0.2
L1 N3 2 18.77u
.ends 4025_74404043220A_22u
*******
.subckt 4025_74404043330A_33u 1 2
Rp 1 2 36000
Cp 1 2 2.18p
Rs 1 N3 0.316
L1 N3 2 29.3u
.ends 4025_74404043330A_33u
*******
.subckt 4025_74404043470A_47u 1 2
Rp 1 2 47600
Cp 1 2 2.3p
Rs 1 N3 0.492
L1 N3 2 39.9u
.ends 4025_74404043470A_47u
*******
.subckt 4025_74404043221A_220u  1 2
Rp 1 2 164796
Cp 1 2 2.493p
Rs 1 N3 2.43
L1 N3 2 200.311u
.ends 4025_74404043221A_220u 
*******
.subckt 4025_74404043471A_470u  1 2
Rp 1 2 992355
Cp 1 2 2.412p
Rs 1 N3 3.55
L1 N3 2 420.135u
.ends 4025_74404043471A_470u 
*******
.subckt 5020_74404052010_1u 1 2
Rp 1 2 2057
Cp 1 2 1.915p
Rs 1 N3 0.0198
L1 N3 2 0.777053u
.ends 5020_74404052010_1u
*******
.subckt 5020_74404052012_1.2u 1 2
Rp 1 2 2139
Cp 1 2 1.407p
Rs 1 N3 0.0234
L1 N3 2 0.989227u
.ends 5020_74404052012_1.2u
*******
.subckt 5020_74404052015_1.5u 1 2
Rp 1 2 3078
Cp 1 2 2.077p
Rs 1 N3 0.0257
L1 N3 2 1.277u
.ends 5020_74404052015_1.5u
*******
.subckt 5020_74404052022_2.2u 1 2
Rp 1 2 3683
Cp 1 2 2.093p
Rs 1 N3 0.0316
L1 N3 2 1.581u
.ends 5020_74404052022_2.2u
*******
.subckt 5020_74404052033_3.3u 1 2
Rp 1 2 5197
Cp 1 2 1.992p
Rs 1 N3 0.0422
L1 N3 2 3.197u
.ends 5020_74404052033_3.3u
*******
.subckt 5020_74404052039_3.9u 1 2
Rp 1 2 4725
Cp 1 2 2.34p
Rs 1 N3 0.0505
L1 N3 2 2.743u
.ends 5020_74404052039_3.9u
*******
.subckt 5020_74404052047_4.7u 1 2
Rp 1 2 6463
Cp 1 2 2.223p
Rs 1 N3 0.0559
L1 N3 2 4.058u
.ends 5020_74404052047_4.7u
*******
.subckt 5020_74404052056_5.6u 1 2
Rp 1 2 6630
Cp 1 2 1.789p
Rs 1 N3 0.0675
L1 N3 2 5.682u
.ends 5020_74404052056_5.6u
*******
.subckt 5020_74404052075_7.5u 1 2
Rp 1 2 9937
Cp 1 2 2.076p
Rs 1 N3 0.0968
L1 N3 2 7.819u
.ends 5020_74404052075_7.5u
*******
.subckt 5020_74404052100_10u 1 2
Rp 1 2 11300
Cp 1 2 2.136p
Rs 1 N3 0.109
L1 N3 2 8.543u
.ends 5020_74404052100_10u
*******
.subckt 5020_74404052101_100u 1 2
Rp 1 2 39059
Cp 1 2 3.805p
Rs 1 N3 1.09
L1 N3 2 89.236u
.ends 5020_74404052101_100u
*******
.subckt 5020_74404052150_15u 1 2
Rp 1 2 14175
Cp 1 2 2.244p
Rs 1 N3 0.162
L1 N3 2 13.122u
.ends 5020_74404052150_15u
*******
.subckt 5020_74404052220_22u 1 2
Rp 1 2 15930
Cp 1 2 3.01p
Rs 1 N3 0.225
L1 N3 2 16.452u
.ends 5020_74404052220_22u
*******
.subckt 5020_74404052330_33u 1 2
Rp 1 2 20038
Cp 1 2 2.925p
Rs 1 N3 0.387
L1 N3 2 32.071u
.ends 5020_74404052330_33u
*******
.subckt 5020_74404052470_47u 1 2
Rp 1 2 20644
Cp 1 2 5.425p
Rs 1 N3 0.521
L1 N3 2 35.145u
.ends 5020_74404052470_47u
*******
.subckt 5020_74404052560_56u 1 2
Rp 1 2 34622
Cp 1 2 2.286p
Rs 1 N3 0.627
L1 N3 2 52.706u
.ends 5020_74404052560_56u
*******
.subckt 5020_74404052680_68u 1 2
Rp 1 2 32847
Cp 1 2 3.513p
Rs 1 N3 0.769
L1 N3 2 64.039u
.ends 5020_74404052680_68u
*******
.subckt 5020_744040520047_0.47u 1 2
Rp 1 2 931.686
Cp 1 2 0.768756p
Rs 1 N3 0.0139
L1 N3 2 0.396143u
.ends 5020_744040520047_0.47u
*******
.subckt 5020_74404052068_6.8u  1 2
Rp 1 2 3076
Cp 1 2 7.38p
Rs 1 N3 0.0827
L1 N3 2 6.8u
.ends 5020_74404052068_6.8u 
*******
.subckt 5040_74404054151_150u 1 2
Rp 1 2 60234
Cp 1 2 4.81p
Rs 1 N3 0.81
L1 N3 2 142.27u
.ends 5040_74404054151_150u
*******
.subckt 5040_74404054221_220u 1 2
Rp 1 2 70590
Cp 1 2 5.38p
Rs 1 N3 1.4
L1 N3 2 228.36u
.ends 5040_74404054221_220u
*******
.subckt 5040_74404054331_330u 1 2
Rp 1 2 87414
Cp 1 2 5.79p
Rs 1 N3 2.1
L1 N3 2 338.88u
.ends 5040_74404054331_330u
*******
.subckt 5040_74404054471_470u 1 2
Rp 1 2 81435
Cp 1 2 9.5p
Rs 1 N3 2.95
L1 N3 2 421.19u
.ends 5040_74404054471_470u
*******
.subckt 5040_74404054681_680u 1 2
Rp 1 2 137682
Cp 1 2 6.422p
Rs 1 N3 3.98
L1 N3 2 692.898u
.ends 5040_74404054681_680u
*******
.subckt 5040_74404054010_1u 1 2
Rp 1 2 2341
Cp 1 2 0.998p
Rs 1 N3 0.012
L1 N3 2 0.802u
.ends 5040_74404054010_1u
*******
.subckt 5040_74404054015_1.5u 1 2
Rp 1 2 3157
Cp 1 2 2.007p
Rs 1 N3 0.015
L1 N3 2 1.399u
.ends 5040_74404054015_1.5u
*******
.subckt 5040_74404054022_2.2u 1 2
Rp 1 2 3747
Cp 1 2 3.2p
Rs 1 N3 0.019
L1 N3 2 1.951u
.ends 5040_74404054022_2.2u
*******
.subckt 5040_74404054033_3.3u 1 2
Rp 1 2 4776
Cp 1 2 3.865p
Rs 1 N3 0.024
L1 N3 2 2.957u
.ends 5040_74404054033_3.3u
*******
.subckt 5040_74404054047_4.7u 1 2
Rp 1 2 6726
Cp 1 2 4.212p
Rs 1 N3 0.03
L1 N3 2 4.161u
.ends 5040_74404054047_4.7u
*******
.subckt 5040_74404054068_6.8u 1 2
Rp 1 2 7484
Cp 1 2 4.835p
Rs 1 N3 0.043
L1 N3 2 5.737u
.ends 5040_74404054068_6.8u
*******
.subckt 5040_74404054100_10u 1 2
Rp 1 2 9907
Cp 1 2 3.988p
Rs 1 N3 0.064
L1 N3 2 9.227u
.ends 5040_74404054100_10u
*******
.subckt 5040_74404054101_100u 1 2
Rp 1 2 39666
Cp 1 2 4.6p
Rs 1 N3 0.56
L1 N3 2 93.13u
.ends 5040_74404054101_100u
*******
.subckt 5040_74404054102_1000u 1 2
Rp 1 2 171858
Cp 1 2 6.722p
Rs 1 N3 6
L1 N3 2 1057u
.ends 5040_74404054102_1000u
*******
.subckt 5040_74404054150_15u 1 2
Rp 1 2 15117
Cp 1 2 4.799p
Rs 1 N3 0.086
L1 N3 2 13.75u
.ends 5040_74404054150_15u
*******
.subckt 5040_74404054220_22u 1 2
Rp 1 2 17030
Cp 1 2 4.96p
Rs 1 N3 0.129
L1 N3 2 18.3u
.ends 5040_74404054220_22u
*******
.subckt 5040_74404054330_33u 1 2
Rp 1 2 19899
Cp 1 2 4.987p
Rs 1 N3 0.188
L1 N3 2 30.028u
.ends 5040_74404054330_33u
*******
.subckt 5040_74404054470_47u 1 2
Rp 1 2 28181
Cp 1 2 6.194p
Rs 1 N3 0.272
L1 N3 2 39.83u
.ends 5040_74404054470_47u
*******
.subckt 5040_74404054680_68u 1 2
Rp 1 2 39993
Cp 1 2 6.05p
Rs 1 N3 0.4
L1 N3 2 64.82u
.ends 5040_74404054680_68u
*******
.subckt 6028_74404063010_1u 1 2
Rp 1 2 1687
Cp 1 2 1.938p
Rs 1 N3 0.01
L1 N3 2 0.883u
.ends 6028_74404063010_1u
*******
.subckt 6028_74404063012_1.2u 1 2
Rp 1 2 2309
Cp 1 2 2.72p
Rs 1 N3 0.012
L1 N3 2 1.036u
.ends 6028_74404063012_1.2u
*******
.subckt 6028_74404063015_1.5u 1 2
Rp 1 2 2358
Cp 1 2 2.252p
Rs 1 N3 0.013
L1 N3 2 1.32u
.ends 6028_74404063015_1.5u
*******
.subckt 6028_74404063022_2.2u 1 2
Rp 1 2 4062
Cp 1 2 2.36p
Rs 1 N3 0.02
L1 N3 2 2.1u
.ends 6028_74404063022_2.2u
*******
.subckt 6028_74404063033_3.3u 1 2
Rp 1 2 5178
Cp 1 2 3.133p
Rs 1 N3 0.025
L1 N3 2 2.77u
.ends 6028_74404063033_3.3u
*******
.subckt 6028_74404063047_4.7u 1 2
Rp 1 2 5518
Cp 1 2 2.868p
Rs 1 N3 0.03
L1 N3 2 4.264u
.ends 6028_74404063047_4.7u
*******
.subckt 6028_74404063068_6.8u 1 2
Rp 1 2 8308
Cp 1 2 2.836p
Rs 1 N3 0.047
L1 N3 2 6.486u
.ends 6028_74404063068_6.8u
*******
.subckt 6028_74404063082_8.2u 1 2
Rp 1 2 8968
Cp 1 2 2.776p
Rs 1 N3 0.055
L1 N3 2 8.303u
.ends 6028_74404063082_8.2u
*******
.subckt 6028_74404063100_10u 1 2
Rp 1 2 10363
Cp 1 2 3.774p
Rs 1 N3 0.072
L1 N3 2 8.046u
.ends 6028_74404063100_10u
*******
.subckt 6028_74404063101_100u 1 2
Rp 1 2 41364
Cp 1 2 4.844p
Rs 1 N3 0.5
L1 N3 2 92.64u
.ends 6028_74404063101_100u
*******
.subckt 6028_74404063102_1000u 1 2
Rp 1 2 220630
Cp 1 2 4.496p
Rs 1 N3 6.44
L1 N3 2 950.95u
.ends 6028_74404063102_1000u
*******
.subckt 6028_74404063150_15u 1 2
Rp 1 2 14108
Cp 1 2 4.077p
Rs 1 N3 0.125
L1 N3 2 13.938u
.ends 6028_74404063150_15u
*******
.subckt 6028_74404063220_22u 1 2
Rp 1 2 15943
Cp 1 2 3.48p
Rs 1 N3 0.14
L1 N3 2 21.33u
.ends 6028_74404063220_22u
*******
.subckt 6028_74404063330_33u 1 2
Rp 1 2 27088
Cp 1 2 3.032p
Rs 1 N3 0.185
L1 N3 2 29.95u
.ends 6028_74404063330_33u
*******
.subckt 6028_74404063470_47u 1 2
Rp 1 2 26057
Cp 1 2 4.057p
Rs 1 N3 0.315
L1 N3 2 41.012u
.ends 6028_74404063470_47u
*******
.subckt 6028_74404063680_68u 1 2
Rp 1 2 37723
Cp 1 2 3.358p
Rs 1 N3 0.36
L1 N3 2 58.33u
.ends 6028_74404063680_68u
*******
.subckt 6028_744040630082_0.82u 1 2
Rp 1 2 1681
Cp 1 2 2.261p
Rs 1 N3 0.01
L1 N3 2 0.69u
.ends 6028_744040630082_0.82u
*******
.subckt 6028_74404063681_680u  1 2
Rp 1 2 372702
Cp 1 2 4.61p
Rs 1 N3 5.526
L1 N3 2 723.317u
.ends 6028_74404063681_680u 
*******
.subckt 6045_74404064331_330u 1 2
Rp 1 2 89667
Cp 1 2 6.424p
Rs 1 N3 1.177
L1 N3 2 305.495u
.ends 6045_74404064331_330u
*******
.subckt 6045_74404064681_680u 1 2
Rp 1 2 105004
Cp 1 2 7.559p
Rs 1 N3 2.65
L1 N3 2 542.013u
.ends 6045_74404064681_680u
*******
.subckt 6045_74404064010_1u 1 2
Rp 1 2 2277
Cp 1 2 1.332p
Rs 1 N3 0.011
L1 N3 2 0.729u
.ends 6045_74404064010_1u
*******
.subckt 6045_74404064015_1.5u 1 2
Rp 1 2 3391
Cp 1 2 2.738p
Rs 1 N3 0.012
L1 N3 2 1.457u
.ends 6045_74404064015_1.5u
*******
.subckt 6045_74404064018_1.8u 1 2
Rp 1 2 3378
Cp 1 2 2.617p
Rs 1 N3 0.012
L1 N3 2 1.528u
.ends 6045_74404064018_1.8u
*******
.subckt 6045_74404064022_2.2u 1 2
Rp 1 2 3376
Cp 1 2 4.642p
Rs 1 N3 0.014
L1 N3 2 1.948u
.ends 6045_74404064022_2.2u
*******
.subckt 6045_74404064033_3.3u 1 2
Rp 1 2 5613
Cp 1 2 5.253p
Rs 1 N3 0.021
L1 N3 2 3.089u
.ends 6045_74404064033_3.3u
*******
.subckt 6045_74404064047_4.7u 1 2
Rp 1 2 7093
Cp 1 2 5.254p
Rs 1 N3 0.026
L1 N3 2 4.388u
.ends 6045_74404064047_4.7u
*******
.subckt 6045_74404064068_6.8u 1 2
Rp 1 2 6893
Cp 1 2 5.251p
Rs 1 N3 0.031
L1 N3 2 5.546u
.ends 6045_74404064068_6.8u
*******
.subckt 6045_74404064082_8.2u 1 2
Rp 1 2 10052
Cp 1 2 5.358p
Rs 1 N3 0.043
L1 N3 2 7.72u
.ends 6045_74404064082_8.2u
*******
.subckt 6045_74404064100_10u 1 2
Rp 1 2 10150
Cp 1 2 7.115p
Rs 1 N3 0.048
L1 N3 2 9.282u
.ends 6045_74404064100_10u
*******
.subckt 6045_74404064101_100u 1 2
Rp 1 2 36787
Cp 1 2 7.954p
Rs 1 N3 0.433
L1 N3 2 86.112u
.ends 6045_74404064101_100u
*******
.subckt 6045_74404064102_1000u 1 2
Rp 1 2 124743
Cp 1 2 7.902p
Rs 1 N3 4.783
L1 N3 2 806.282u
.ends 6045_74404064102_1000u
*******
.subckt 6045_74404064120_12u 1 2
Rp 1 2 9899
Cp 1 2 7.566p
Rs 1 N3 0.058
L1 N3 2 9.065u
.ends 6045_74404064120_12u
*******
.subckt 6045_74404064121_120u 1 2
Rp 1 2 49057
Cp 1 2 7.21p
Rs 1 N3 0.52
L1 N3 2 93.103u
.ends 6045_74404064121_120u
*******
.subckt 6045_74404064150_15u 1 2
Rp 1 2 13652
Cp 1 2 7.041p
Rs 1 N3 0.068
L1 N3 2 13.321u
.ends 6045_74404064150_15u
*******
.subckt 6045_74404064151_150u 1 2
Rp 1 2 49043
Cp 1 2 6.191p
Rs 1 N3 0.57
L1 N3 2 116.571u
.ends 6045_74404064151_150u
*******
.subckt 6045_74404064180_18u 1 2
Rp 1 2 12232
Cp 1 2 6.707p
Rs 1 N3 0.081
L1 N3 2 13.984u
.ends 6045_74404064180_18u
*******
.subckt 6045_74404064220_22u 1 2
Rp 1 2 15329
Cp 1 2 6.385p
Rs 1 N3 0.089
L1 N3 2 20.865u
.ends 6045_74404064220_22u
*******
.subckt 6045_74404064221_220u 1 2
Rp 1 2 67135
Cp 1 2 6.695p
Rs 1 N3 0.85
L1 N3 2 206.373u
.ends 6045_74404064221_220u
*******
.subckt 6045_74404064330_33u 1 2
Rp 1 2 23074
Cp 1 2 6.43p
Rs 1 N3 0.137
L1 N3 2 29.425u
.ends 6045_74404064330_33u
*******
.subckt 6045_74404064470_47u 1 2
Rp 1 2 23991
Cp 1 2 7.089p
Rs 1 N3 0.2
L1 N3 2 42.609u
.ends 6045_74404064470_47u
*******
.subckt 6045_74404064560_56u 1 2
Rp 1 2 20957
Cp 1 2 9.372p
Rs 1 N3 0.22
L1 N3 2 41.15u
.ends 6045_74404064560_56u
*******
.subckt 6045_74404064680_68u 1 2
Rp 1 2 33997
Cp 1 2 6.624p
Rs 1 N3 0.289
L1 N3 2 64.775u
.ends 6045_74404064680_68u
*******
.subckt 6045_74404064012_1.2u  1 2
Rp 1 2 2842.9
Cp 1 2 1.65126p
Rs 1 N3 0.01
L1 N3 2 1.2u
.ends 6045_74404064012_1.2u 
*******
.subckt 6045_744040640047_0.47u  1 2
Rp 1 2 1691
Cp 1 2 1.091p
Rs 1 N3 0.006
L1 N3 2 0.47u
.ends 6045_744040640047_0.47u 
*******
.subckt 6045_744040640068_0.68u  1 2
Rp 1 2 1552
Cp 1 2 1.595p
Rs 1 N3 0.01
L1 N3 2 0.68u
.ends 6045_744040640068_0.68u 
*******
.subckt 8040_74404084010_1u 1 2
Rp 1 2 1984
Cp 1 2 2.3p
Rs 1 N3 0.008
L1 N3 2 0.898u
.ends 8040_74404084010_1u
*******
.subckt 8040_74404084015_1.5u 1 2
Rp 1 2 3200
Cp 1 2 2.3p
Rs 1 N3 0.01
L1 N3 2 1.36u
.ends 8040_74404084015_1.5u
*******
.subckt 8040_74404084022_2.2u 1 2
Rp 1 2 3750
Cp 1 2 4.1p
Rs 1 N3 0.012
L1 N3 2 1.8u
.ends 8040_74404084022_2.2u
*******
.subckt 8040_74404084033_3.3u 1 2
Rp 1 2 5080
Cp 1 2 4.76p
Rs 1 N3 0.017
L1 N3 2 3.41u
.ends 8040_74404084033_3.3u
*******
.subckt 8040_74404084047_4.7u 1 2
Rp 1 2 6850
Cp 1 2 5.7p
Rs 1 N3 0.019
L1 N3 2 4.5u
.ends 8040_74404084047_4.7u
*******
.subckt 8040_74404084068_6.8u 1 2
Rp 1 2 9480
Cp 1 2 5.6p
Rs 1 N3 0.024
L1 N3 2 6.2u
.ends 8040_74404084068_6.8u
*******
.subckt 8040_74404084082_8.2u 1 2
Rp 1 2 9210
Cp 1 2 5.6p
Rs 1 N3 0.026
L1 N3 2 8.18u
.ends 8040_74404084082_8.2u
*******
.subckt 8040_74404084100_10u 1 2
Rp 1 2 11920
Cp 1 2 5.3p
Rs 1 N3 0.029
L1 N3 2 8.7u
.ends 8040_74404084100_10u
*******
.subckt 8040_74404084101_100u 1 2
Rp 1 2 36750
Cp 1 2 8.3p
Rs 1 N3 0.29
L1 N3 2 92.2u
.ends 8040_74404084101_100u
*******
.subckt 8040_74404084102_1000u 1 2
Rp 1 2 167100
Cp 1 2 5.79p
Rs 1 N3 2.87
L1 N3 2 970.7u
.ends 8040_74404084102_1000u
*******
.subckt 8040_74404084120_12u 1 2
Rp 1 2 15750
Cp 1 2 5.56p
Rs 1 N3 0.04
L1 N3 2 10.2u
.ends 8040_74404084120_12u
*******
.subckt 8040_74404084121_120u 1 2
Rp 1 2 42120
Cp 1 2 6.7p
Rs 1 N3 0.347
L1 N3 2 113.2u
.ends 8040_74404084121_120u
*******
.subckt 8040_74404084150_15u 1 2
Rp 1 2 11370
Cp 1 2 6.9p
Rs 1 N3 0.047
L1 N3 2 15.18u
.ends 8040_74404084150_15u
*******
.subckt 8040_74404084151_150u 1 2
Rp 1 2 40102
Cp 1 2 8.651p
Rs 1 N3 0.478
L1 N3 2 118.98u
.ends 8040_74404084151_150u
*******
.subckt 8040_74404084180_18u 1 2
Rp 1 2 19840
Cp 1 2 6.4p
Rs 1 N3 0.053
L1 N3 2 14.7u
.ends 8040_74404084180_18u
*******
.subckt 8040_74404084220_22u 1 2
Rp 1 2 20200
Cp 1 2 5.4p
Rs 1 N3 0.069
L1 N3 2 18.9u
.ends 8040_74404084220_22u
*******
.subckt 8040_74404084221_220u 1 2
Rp 1 2 48204
Cp 1 2 8.754p
Rs 1 N3 0.592
L1 N3 2 161.599u
.ends 8040_74404084221_220u
*******
.subckt 8040_74404084330_33u 1 2
Rp 1 2 19670
Cp 1 2 7p
Rs 1 N3 0.097
L1 N3 2 30.1u
.ends 8040_74404084330_33u
*******
.subckt 8040_74404084331_330u 1 2
Rp 1 2 74300
Cp 1 2 7.4p
Rs 1 N3 0.865
L1 N3 2 296.5u
.ends 8040_74404084331_330u
*******
.subckt 8040_74404084470_47u 1 2
Rp 1 2 22230
Cp 1 2 9.1p
Rs 1 N3 0.136
L1 N3 2 44.7u
.ends 8040_74404084470_47u
*******
.subckt 8040_74404084560_56u 1 2
Rp 1 2 27870
Cp 1 2 7.9p
Rs 1 N3 0.18
L1 N3 2 51.4u
.ends 8040_74404084560_56u
*******
.subckt 8040_74404084680_68u 1 2
Rp 1 2 29330
Cp 1 2 7.8p
Rs 1 N3 0.196
L1 N3 2 61.8u
.ends 8040_74404084680_68u
*******
.subckt 8040_74404084681_680u 1 2
Rp 1 2 122365
Cp 1 2 6.864p
Rs 1 N3 2.032
L1 N3 2 630.57u
.ends 8040_74404084681_680u
*******
.subckt 8065_74404086221_220u 1 2
Rp 1 2 59302
Cp 1 2 15.439p
Rs 1 N3 0.555
L1 N3 2 190.032u
.ends 8065_74404086221_220u
*******
.subckt 8065_74404086102_1000u 1 2
Rp 1 2 120450
Cp 1 2 11.668p
Rs 1 N3 2.35
L1 N3 2 864.742u
.ends 8065_74404086102_1000u
*******
.subckt 8065_74404086152_1500u 1 2
Rp 1 2 137739
Cp 1 2 15.7690877865p
Rs 1 N3 3.65
L1 N3 2 1428.972772943u
.ends 8065_74404086152_1500u
*******
.subckt 8065_74404086222_2200u 1 2
Rp 1 2 227946
Cp 1 2 15.81587720877p
Rs 1 N3 5
L1 N3 2 1947.832355291u
.ends 8065_74404086222_2200u
*******
.subckt 8065_74404086332_3300u 1 2
Rp 1 2 267101
Cp 1 2 10.386p
Rs 1 N3 7.3
L1 N3 2 3128u
.ends 8065_74404086332_3300u
*******
.subckt 8065_74404086472_4700u 1 2
Rp 1 2 295575
Cp 1 2 13.635p
Rs 1 N3 12.15
L1 N3 2 4277u
.ends 8065_74404086472_4700u
*******
.subckt 8065_74404086682_6800u 1 2
Rp 1 2 371955
Cp 1 2 13.058p
Rs 1 N3 18.7
L1 N3 2 6342u
.ends 8065_74404086682_6800u
*******
.subckt 8065_74404086101_100u  1 2
Rp 1 2 49550
Cp 1 2 15.52p
Rs 1 N3 0.238
L1 N3 2 94.56u
.ends 8065_74404086101_100u 
*******
.subckt 8065_74404086103_10000u  1 2
Rp 1 2 443000
Cp 1 2 17.65p
Rs 1 N3 22.8
L1 N3 2 8836u
.ends 8065_74404086103_10000u 
*******
.subckt 8065_74404086151_150u  1 2
Rp 1 2 66107
Cp 1 2 15.97p
Rs 1 N3 0.355
L1 N3 2 139.75u
.ends 8065_74404086151_150u 
*******
.subckt 8065_74404086331_330u  1 2
Rp 1 2 93840
Cp 1 2 14.79p
Rs 1 N3 0.7
L1 N3 2 310.97u
.ends 8065_74404086331_330u 
*******
.subckt 8065_74404086471_470u  1 2
Rp 1 2 106610
Cp 1 2 16.92p
Rs 1 N3 1.2
L1 N3 2 493.31u
.ends 8065_74404086471_470u 
*******
.subckt 8065_74404086681_680u  1 2
Rp 1 2 109785
Cp 1 2 14.707p
Rs 1 N3 1.65
L1 N3 2 651.45u
.ends 8065_74404086681_680u 
*******
