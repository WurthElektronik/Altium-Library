**************************************************
* Manufacturer:          Würth Elektronik 
* Kinds:                 Multilayer Ceramic Chip Capacitors
* Matchcode:             WCAP-CSSA
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1808_8853520100071_33pF 1 2
Rser 1 3 0.131840103427
Lser 2 4 0.00000000095
C1 3 4 0.000000000033
Rpar 3 4 100000000000
.ends 1808_8853520100071_33pF
*******
.subckt 1808_8853522100131_1nF 1 2
Rser 1 3 0.19143371088
Lser 2 4 0.0000000008
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1808_8853522100131_1nF
*******
.subckt 1812_8853522110011_470pF 1 2
Rser 1 3 0.235
Lser 2 4 0.000000000505
C1 3 4 0.00000000047
Rpar 3 4 100000000000
.ends 1812_8853522110011_470pF
*******
.subckt 1812_8853522110021_680pF 1 2
Rser 1 3 0.192401658822
Lser 2 4 0.0000000005
C1 3 4 0.00000000068
Rpar 3 4 100000000000
.ends 1812_8853522110021_680pF
*******
.subckt 1812_8853522110031_1nF 1 2
Rser 1 3 0.17
Lser 2 4 0.00000000081
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_8853522110031_1nF
*******
.subckt 2211_8853522130111_1nF 1 2
Rser 1 3 0.15
Lser 2 4 1.080985281E-09
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 2211_8853522130111_1nF
*******
.subckt 2211_8853522130151_2.2nF 1 2
Rser 1 3 0.1
Lser 2 4 1.052883757E-09
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 2211_8853522130151_2.2nF
*******
.subckt 2220_8853522140011_4.7nF 1 2
Rser 1 3 0.0355
Lser 2 4 0.0000000005
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 2220_8853522140011_4.7nF
*******
.subckt 1808_8853620100091_33pF 1 2
Rser 1 3 0.35
Lser 2 4 0.00000000075
C1 3 4 0.000000000033
Rpar 3 4 100000000000
.ends 1808_8853620100091_33pF
*******
.subckt 1808_8853620100111_47pF 1 2
Rser 1 3 0.16
Lser 2 4 0.000000001
C1 3 4 0.000000000047
Rpar 3 4 100000000000
.ends 1808_8853620100111_47pF
*******
.subckt 1808_8853620100171_100pF 1 2
Rser 1 3 0.0287431979621
Lser 2 4 0.0000000011
C1 3 4 0.0000000001
Rpar 3 4 100000000000
.ends 1808_8853620100171_100pF
*******
.subckt 1808_8853620100181_220pF 1 2
Rser 1 3 0.0587493769172
Lser 2 4 0.00000000095
C1 3 4 0.00000000022
Rpar 3 4 100000000000
.ends 1808_8853620100181_220pF
*******
.subckt 1808_8853622100091_470pF 1 2
Rser 1 3 0.27
Lser 2 4 0.00000000066
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1808_8853622100091_470pF
*******
.subckt 1808_8853622100131_680pF 1 2
Rser 1 3 0.19
Lser 2 4 7.08923866E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1808_8853622100131_680pF
*******
.subckt 1808_8853622100171_1nF 1 2
Rser 1 3 0.215
Lser 2 4 0.00000000075
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1808_8853622100171_1nF
*******
.subckt 1808_8853622100181_150pF 1 2
Rser 1 3 0.48
Lser 2 4 0.000000000615
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1808_8853622100181_150pF
*******
.subckt 1812_8853622110111_1nF 1 2
Rser 1 3 0.15
Lser 2 4 5.98981061E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_8853622110111_1nF
*******
.subckt 1812_8853622110151_2.2nF 1 2
Rser 1 3 0.120953454829
Lser 2 4 8.07194919E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1812_8853622110151_2.2nF
*******
