**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Power Multilayer Inductor
* Matchcode:              WE-PMI 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1008_74479787147B_0.47u 1 2
Rp 1 2 600
Cp 1 2 4.1p
Rs 1 N3 0.04
L1 N3 2 0.47u
.ends 1008_74479787147B_0.47u
*******
.subckt 1008_74479787210B_1u 1 2
Rp 1 2 1100
Cp 1 2 4p
Rs 1 N3 0.06
L1 N3 2 1u
.ends 1008_74479787210B_1u
*******
.subckt 1008_74479787215A_1.5u 1 2
Rp 1 2 1650
Cp 1 2 3.8p
Rs 1 N3 0.07
L1 N3 2 1.5u
.ends 1008_74479787215A_1.5u
*******
.subckt 1008_74479787222A_2.2u 1 2
Rp 1 2 2100
Cp 1 2 3.6p
Rs 1 N3 0.085
L1 N3 2 2.2u
.ends 1008_74479787222A_2.2u
*******
.subckt 1008_74479787233A_3.3u 1 2
Rp 1 2 2100
Cp 1 2 3.5p
Rs 1 N3 0.1
L1 N3 2 3.3u
.ends 1008_74479787233A_3.3u
*******
.subckt 1008_74479787247A_4.7u 1 2
Rp 1 2 2200
Cp 1 2 3.5p
Rs 1 N3 0.11
L1 N3 2 4.7u
.ends 1008_74479787247A_4.7u
*******
.subckt 1008_74479887124C_0.24u 1 2
Rp 1 2 525.038
Cp 1 2 4.02p
Rs 1 N3 0.02
L1 N3 2 0.24u
.ends 1008_74479887124C_0.24u
*******
.subckt 1008_74479887147C_0.47u 1 2
Rp 1 2 1031.41
Cp 1 2 3.567p
Rs 1 N3 0.033
L1 N3 2 0.47u
.ends 1008_74479887147C_0.47u
*******
.subckt 1008_74479887210C_1u 1 2
Rp 1 2 1564.25
Cp 1 2 4.613p
Rs 1 N3 0.045
L1 N3 2 1u
.ends 1008_74479887210C_1u
*******
.subckt 1008_74479887222C_2.2u 1 2
Rp 1 2 2962.14
Cp 1 2 2.929p
Rs 1 N3 0.09
L1 N3 2 2.2u
.ends 1008_74479887222C_2.2u
*******
.subckt 1008_74479889268_6.8u 1 2
Rp 1 2 7000
Cp 1 2 2.8p
Rs 1 N3 0.5
L1 N3 2 6.8u
.ends 1008_74479889268_6.8u
*******
.subckt 1210_74479897122_0.22u 1 2
Rp 1 2 288.07
Cp 1 2 3.69p
Rs 1 N3 0.016
L1 N3 2 0.22u
.ends 1210_74479897122_0.22u
*******
.subckt 1210_74479897150_0.5u 1 2
Rp 1 2 466.11
Cp 1 2 3.731p
Rs 1 N3 0.025
L1 N3 2 0.5u
.ends 1210_74479897150_0.5u
*******
.subckt 1210_74479899111_0.11u 1 2
Rp 1 2 166.683
Cp 1 2 2.105p
Rs 1 N3 0.007
L1 N3 2 0.11u
.ends 1210_74479899111_0.11u
*******
.subckt 1210_74479899130_0.3u 1 2
Rp 1 2 362.407
Cp 1 2 4.338p
Rs 1 N3 0.015
L1 N3 2 0.3u
.ends 1210_74479899130_0.3u
*******
.subckt 1210_74479899150_0.5u 1 2
Rp 1 2 641.519
Cp 1 2 3.012p
Rs 1 N3 0.018
L1 N3 2 0.5u
.ends 1210_74479899150_0.5u
*******
.subckt 1210_74479899210_1u 1 2
Rp 1 2 1469
Cp 1 2 3.439p
Rs 1 N3 0.05
L1 N3 2 1u
.ends 1210_74479899210_1u
*******
.subckt 0603_74479762122_0.22u 1 2
Rp 1 2 600
Cp 1 2 1.4p
Rs 1 N3 0.12
L1 N3 2 0.22u
.ends 0603_74479762122_0.22u
*******
.subckt 0603_74479762133_0.33u 1 2
Rp 1 2 850
Cp 1 2 1.55p
Rs 1 N3 0.16
L1 N3 2 0.33u
.ends 0603_74479762133_0.33u
*******
.subckt 0603_74479762168_0.68u 1 2
Rp 1 2 1200
Cp 1 2 1.4p
Rs 1 N3 0.22
L1 N3 2 0.68u
.ends 0603_74479762168_0.68u
*******
.subckt 0603_74479763147_0.47u 1 2
Rp 1 2 600
Cp 1 2 1.1p
Rs 1 N3 0.3
L1 N3 2 0.47u
.ends 0603_74479763147_0.47u
*******
.subckt 0603_74479763147A_0.47u 1 2
Rp 1 2 1200
Cp 1 2 1.45p
Rs 1 N3 0.09
L1 N3 2 0.47u
.ends 0603_74479763147A_0.47u
*******
.subckt 0603_74479763168_0.68u 1 2
Rp 1 2 1500
Cp 1 2 1.2p
Rs 1 N3 0.18
L1 N3 2 0.68u
.ends 0603_74479763168_0.68u
*******
.subckt 0603_74479763210_1u 1 2
Rp 1 2 1000
Cp 1 2 1.1p
Rs 1 N3 0.3
L1 N3 2 1u
.ends 0603_74479763210_1u
*******
.subckt 0603_74479763210A_1u 1 2
Rp 1 2 1600
Cp 1 2 1.25p
Rs 1 N3 0.2
L1 N3 2 1u
.ends 0603_74479763210A_1u
*******
.subckt 0603_74479763215_1.5u 1 2
Rp 1 2 2000
Cp 1 2 1.3p
Rs 1 N3 0.23
L1 N3 2 1.5u
.ends 0603_74479763215_1.5u
*******
.subckt 0603_74479763222_2.2u 1 2
Rp 1 2 2100
Cp 1 2 1.35p
Rs 1 N3 0.3
L1 N3 2 2.2u
.ends 0603_74479763222_2.2u
*******
.subckt 0805_74479773133_0.33u 1 2
Rp 1 2 650
Cp 1 2 2p
Rs 1 N3 0.1
L1 N3 2 0.33u
.ends 0805_74479773133_0.33u
*******
.subckt 0805_74479773147_0.47u 1 2
Rp 1 2 900
Cp 1 2 2.2p
Rs 1 N3 0.1
L1 N3 2 0.47u
.ends 0805_74479773147_0.47u
*******
.subckt 0805_74479773154_0.54u 1 2
Rp 1 2 920
Cp 1 2 2.2p
Rs 1 N3 0.12
L1 N3 2 0.54u
.ends 0805_74479773154_0.54u
*******
.subckt 0805_74479773210_1u 1 2
Rp 1 2 1600
Cp 1 2 2.2p
Rs 1 N3 0.18
L1 N3 2 1u
.ends 0805_74479773210_1u
*******
.subckt 0805_74479774147_0.47u 1 2
Rp 1 2 550
Cp 1 2 1.75p
Rs 1 N3 0.12
L1 N3 2 0.47u
.ends 0805_74479774147_0.47u
*******
.subckt 0805_74479774210_1u 1 2
Rp 1 2 1200
Cp 1 2 2p
Rs 1 N3 0.19
L1 N3 2 1u
.ends 0805_74479774210_1u
*******
.subckt 0805_74479774215_1.5u 1 2
Rp 1 2 1800
Cp 1 2 1.55p
Rs 1 N3 0.26
L1 N3 2 1.5u
.ends 0805_74479774215_1.5u
*******
.subckt 0805_74479774222_2.2u 1 2
Rp 1 2 2300
Cp 1 2 2.2p
Rs 1 N3 0.34
L1 N3 2 2.2u
.ends 0805_74479774222_2.2u
*******
.subckt 0805_74479775147A_0.47u 1 2
Rp 1 2 1000
Cp 1 2 1.3p
Rs 1 N3 0.1
L1 N3 2 0.47u
.ends 0805_74479775147A_0.47u
*******
.subckt 0805_74479775210A_1u 1 2
Rp 1 2 1600
Cp 1 2 2p
Rs 1 N3 0.11
L1 N3 2 1u
.ends 0805_74479775210A_1u
*******
.subckt 0805_74479775215_1.5u 1 2
Rp 1 2 1800
Cp 1 2 2p
Rs 1 N3 0.16
L1 N3 2 1.5u
.ends 0805_74479775215_1.5u
*******
.subckt 0805_74479775222A_2.2u 1 2
Rp 1 2 2000
Cp 1 2 2.1p
Rs 1 N3 0.2
L1 N3 2 2.2u
.ends 0805_74479775222A_2.2u
*******
.subckt 0805_74479775233_3.3u 1 2
Rp 1 2 2000
Cp 1 2 2.2p
Rs 1 N3 0.2
L1 N3 2 3.3u
.ends 0805_74479775233_3.3u
*******
.subckt 0805_74479775247_4.7u 1 2
Rp 1 2 2700
Cp 1 2 2p
Rs 1 N3 0.25
L1 N3 2 4.7u
.ends 0805_74479775247_4.7u
*******
.subckt 0805_74479777268_6.8u 1 2
Rp 1 2 4000
Cp 1 2 2p
Rs 1 N3 0.3
L1 N3 2 6.8u
.ends 0805_74479777268_6.8u
*******
.subckt 0805_74479777310_10u 1 2
Rp 1 2 9000
Cp 1 2 2.5p
Rs 1 N3 0.5
L1 N3 2 10u
.ends 0805_74479777310_10u
*******
.subckt 0805_74479777310A_10u 1 2
Rp 1 2 4000
Cp 1 2 2.1p
Rs 1 N3 0.3
L1 N3 2 10u
.ends 0805_74479777310A_10u
*******
.subckt 0805_74479875210C_1u 1 2
Rp 1 2 1719.82
Cp 1 2 1.763p
Rs 1 N3 0.115
L1 N3 2 1u
.ends 0805_74479875210C_1u
*******
.subckt 0805_74479875222C_2.2u 1 2
Rp 1 2 2277.85
Cp 1 2 2.151p
Rs 1 N3 0.14
L1 N3 2 2.2u
.ends 0805_74479875222C_2.2u
*******
.subckt 0805LR_74479775147_0.47u 1 2
Rp 1 2 625
Cp 1 2 1.65p
Rs 1 N3 0.075
L1 N3 2 0.47u
.ends 0805LR_74479775147_0.47u
*******
.subckt 0805LR_74479775210_1u 1 2
Rp 1 2 900
Cp 1 2 1.8p
Rs 1 N3 0.1
L1 N3 2 1u
.ends 0805LR_74479775210_1u
*******
.subckt 0805LR_74479775222_2.2u 1 2
Rp 1 2 2300
Cp 1 2 1.8p
Rs 1 N3 0.23
L1 N3 2 2.2u
.ends 0805LR_74479775222_2.2u
*******
.subckt 0806_74479776147_0.47u 1 2
Rp 1 2 1150
Cp 1 2 2.4p
Rs 1 N3 0.08
L1 N3 2 0.47u
.ends 0806_74479776147_0.47u
*******
.subckt 0806_74479776210_1u 1 2
Rp 1 2 1300
Cp 1 2 2.5p
Rs 1 N3 0.09
L1 N3 2 1u
.ends 0806_74479776210_1u
*******
.subckt 0806_74479776215_1.5u 1 2
Rp 1 2 2000
Cp 1 2 2.35p
Rs 1 N3 0.11
L1 N3 2 1.5u
.ends 0806_74479776215_1.5u
*******
.subckt 0806_74479776222A_2.2u 1 2
Rp 1 2 2000
Cp 1 2 2.3p
Rs 1 N3 0.11
L1 N3 2 2.2u
.ends 0806_74479776222A_2.2u
*******
.subckt 0806_74479776233A_3.3u 1 2
Rp 1 2 2100
Cp 1 2 2.3p
Rs 1 N3 0.12
L1 N3 2 3.3u
.ends 0806_74479776233A_3.3u
*******
.subckt 0806_74479776247A_4.7u 1 2
Rp 1 2 2300
Cp 1 2 2.4p
Rs 1 N3 0.14
L1 N3 2 4.7u
.ends 0806_74479776247A_4.7u
*******
.subckt 0806_74479778268_6.8u 1 2
Rp 1 2 3000
Cp 1 2 2p
Rs 1 N3 0.17
L1 N3 2 6.8u
.ends 0806_74479778268_6.8u
*******
.subckt 0806_74479778310_10u 1 2
Rp 1 2 1500
Cp 1 2 2.8p
Rs 1 N3 0.25
L1 N3 2 10u
.ends 0806_74479778310_10u
*******
.subckt 0806_74479876124C_0.24u 1 2
Rp 1 2 395.202
Cp 1 2 8.902p
Rs 1 N3 0.026
L1 N3 2 0.24u
.ends 0806_74479876124C_0.24u
*******
.subckt 0806_74479876147_0.47u 1 2
Rp 1 2 900
Cp 1 2 2.7p
Rs 1 N3 0.04
L1 N3 2 0.47u
.ends 0806_74479876147_0.47u
*******
.subckt 0806_74479876147C_0.47u 1 2
Rp 1 2 652.377
Cp 1 2 9.394p
Rs 1 N3 0.044
L1 N3 2 0.47u
.ends 0806_74479876147C_0.47u
*******
.subckt 0806_74479876168_0.68u 1 2
Rp 1 2 1200
Cp 1 2 3.2p
Rs 1 N3 0.06
L1 N3 2 0.68u
.ends 0806_74479876168_0.68u
*******
.subckt 0806_74479876168C_0.68u 1 2
Rp 1 2 1061.49
Cp 1 2 2.742p
Rs 1 N3 0.068
L1 N3 2 0.68u
.ends 0806_74479876168C_0.68u
*******
.subckt 0806_74479876210_1u 1 2
Rp 1 2 1500
Cp 1 2 2.8p
Rs 1 N3 0.07
L1 N3 2 1u
.ends 0806_74479876210_1u
*******
.subckt 0806_74479876210C_1u 1 2
Rp 1 2 1132.58
Cp 1 2 2.879p
Rs 1 N3 0.075
L1 N3 2 1u
.ends 0806_74479876210C_1u
*******
.subckt 0806_74479876215C_1.5u 1 2
Rp 1 2 2007.8
Cp 1 2 2.147p
Rs 1 N3 0.115
L1 N3 2 1.5u
.ends 0806_74479876215C_1.5u
*******
.subckt 0806_74479876222C_2.2u 1 2
Rp 1 2 3032.39
Cp 1 2 2.285p
Rs 1 N3 0.21
L1 N3 2 2.2u
.ends 0806_74479876222C_2.2u
*******
.subckt 0806HS_74479776222_2.2u 1 2
Rp 1 2 1600
Cp 1 2 1.8p
Rs 1 N3 0.11
L1 N3 2 2.2u
.ends 0806HS_74479776222_2.2u
*******
.subckt 0806HS_74479776233_3.3u 1 2
Rp 1 2 2400
Cp 1 2 1.7p
Rs 1 N3 0.13
L1 N3 2 3.3u
.ends 0806HS_74479776233_3.3u
*******
.subckt 0806HS_74479776247_4.7u 1 2
Rp 1 2 3000
Cp 1 2 1.8p
Rs 1 N3 0.16
L1 N3 2 4.7u
.ends 0806HS_74479776247_4.7u
*******
.subckt 1008_74479888222_2.2u 1 2
Rp 1 2 3600
Cp 1 2 2.6p
Rs 1 N3 0.2
L1 N3 2 2.2u
.ends 1008_74479888222_2.2u
*******
.subckt 1008_74479888233_3.3u 1 2
Rp 1 2 4000
Cp 1 2 2.7p
Rs 1 N3 0.25
L1 N3 2 3.3u
.ends 1008_74479888233_3.3u
*******
.subckt 1008_74479888247_4.7u 1 2
Rp 1 2 5500
Cp 1 2 3.2p
Rs 1 N3 0.38
L1 N3 2 4.7u
.ends 1008_74479888247_4.7u
*******
.subckt 1008_74479888268_6.8u 1 2
Rp 1 2 6500
Cp 1 2 3p
Rs 1 N3 0.45
L1 N3 2 6.8u
.ends 1008_74479888268_6.8u
*******
.subckt 1008_74479888310_10u 1 2
Rp 1 2 6000
Cp 1 2 2.8p
Rs 1 N3 0.5
L1 N3 2 10u
.ends 1008_74479888310_10u
*******
.subckt 1008_74479889210_1u 1 2
Rp 1 2 2400
Cp 1 2 3p
Rs 1 N3 0.085
L1 N3 2 1u
.ends 1008_74479889210_1u
*******
.subckt 1008_74479889222_2.2u 1 2
Rp 1 2 4400
Cp 1 2 2.7p
Rs 1 N3 0.25
L1 N3 2 2.2u
.ends 1008_74479889222_2.2u
*******
.subckt 1008_74479889233_3.3u 1 2
Rp 1 2 6000
Cp 1 2 2.8p
Rs 1 N3 0.25
L1 N3 2 3.3u
.ends 1008_74479889233_3.3u
*******
.subckt 1008_74479889247_4.7u 1 2
Rp 1 2 7500
Cp 1 2 2.8p
Rs 1 N3 0.4
L1 N3 2 4.7u
.ends 1008_74479889247_4.7u
*******
.subckt 1008_74479889310_10u 1 2
Rp 1 2 7800
Cp 1 2 2.9p
Rs 1 N3 0.5
L1 N3 2 10u
.ends 1008_74479889310_10u
*******
.subckt 1008LP_74479787147A_0.47u 1 2
Rp 1 2 300
Cp 1 2 3.1p
Rs 1 N3 0.04
L1 N3 2 0.47u
.ends 1008LP_74479787147A_0.47u
*******
.subckt 1008LP_74479787210A_1u 1 2
Rp 1 2 1000
Cp 1 2 2p
Rs 1 N3 0.055
L1 N3 2 1u
.ends 1008LP_74479787210A_1u
*******
.subckt 1008LP_74479787215_1.5u 1 2
Rp 1 2 1700
Cp 1 2 2.8p
Rs 1 N3 0.07
L1 N3 2 1.5u
.ends 1008LP_74479787215_1.5u
*******
.subckt 1008LP_74479787222_2.2u 1 2
Rp 1 2 2100
Cp 1 2 2.6p
Rs 1 N3 0.08
L1 N3 2 2.2u
.ends 1008LP_74479787222_2.2u
*******
.subckt 1008LP_74479787233_3.3u 1 2
Rp 1 2 2700
Cp 1 2 2.6p
Rs 1 N3 0.1
L1 N3 2 3.3u
.ends 1008LP_74479787233_3.3u
*******
.subckt 1008LP_74479787247_4.7u 1 2
Rp 1 2 3000
Cp 1 2 2.5p
Rs 1 N3 0.11
L1 N3 2 4.7u
.ends 1008LP_74479787247_4.7u
*******
.subckt 1008LP_74479887210A_1u 1 2
Rp 1 2 950
Cp 1 2 2.6p
Rs 1 N3 0.1
L1 N3 2 1u
.ends 1008LP_74479887210A_1u
*******
.subckt 1008LP_74479887222A_2.2u 1 2
Rp 1 2 1400
Cp 1 2 2.3p
Rs 1 N3 0.14
L1 N3 2 2.2u
.ends 1008LP_74479887222A_2.2u
*******
.subckt 1008LP_74479887233A_3.3u 1 2
Rp 1 2 2600
Cp 1 2 2p
Rs 1 N3 0.18
L1 N3 2 3.3u
.ends 1008LP_74479887233A_3.3u
*******
.subckt 1008LP_74479887247A_4.7u 1 2
Rp 1 2 2900
Cp 1 2 2p
Rs 1 N3 0.23
L1 N3 2 4.7u
.ends 1008LP_74479887247A_4.7u
*******
.subckt 1008LP_74479887268A_6.8u 1 2
Rp 1 2 4000
Cp 1 2 1.9p
Rs 1 N3 0.25
L1 N3 2 6.8u
.ends 1008LP_74479887268A_6.8u
*******
.subckt 1008LP_74479887310A_10u 1 2
Rp 1 2 4200
Cp 1 2 1.9p
Rs 1 N3 0.3
L1 N3 2 10u
.ends 1008LP_74479887310A_10u
*******
