**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT High Saturation Power Inductor
* Matchcode:              WE-LQSH
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 2010_744050200047_0.47u 1 2
Rp 1 2 994
Cp 1 2 2.639p
Rs 1 N3 0.041
L1 N3 2 0.47u
.ends 2010_744050200047_0.47u
*******
.subckt 2010_74405020010_1u 1 2
Rp 1 2 1324
Cp 1 2 4.171p
Rs 1 N3 0.075
L1 N3 2 1u
.ends 2010_74405020010_1u
*******
.subckt 2010_74405020015_1.5u 1 2
Rp 1 2 1908
Cp 1 2 3.525p
Rs 1 N3 0.11
L1 N3 2 1.5u
.ends 2010_74405020015_1.5u
*******
.subckt 2010_74405020022_2.5u 1 2
Rp 1 2 2452
Cp 1 2 4.865p
Rs 1 N3 0.142
L1 N3 2 2.5u
.ends 2010_74405020022_2.5u
*******
.subckt 2010_74405020047_4.7u 1 2
Rp 1 2 5078
Cp 1 2 4.451p
Rs 1 N3 0.37
L1 N3 2 4.7u
.ends 2010_74405020047_4.7u
*******
.subckt 2010_74405020100_10u 1 2
Rp 1 2 7894
Cp 1 2 5.459p
Rs 1 N3 0.68
L1 N3 2 10u
.ends 2010_74405020100_10u
*******
.subckt 2512_744050240047_0.47u 1 2
Rp 1 2 777
Cp 1 2 4.138p
Rs 1 N3 0.029
L1 N3 2 0.47u
.ends 2512_744050240047_0.47u
*******
.subckt 2512_74405024010_1u 1 2
Rp 1 2 1145
Cp 1 2 6.529p
Rs 1 N3 0.048
L1 N3 2 1u
.ends 2512_74405024010_1u
*******
.subckt 2512_74405024015_1.5u 1 2
Rp 1 2 1625
Cp 1 2 6.589p
Rs 1 N3 0.06
L1 N3 2 1.5u
.ends 2512_74405024015_1.5u
*******
.subckt 2512_74405024022_2.2u 1 2
Rp 1 2 2054
Cp 1 2 6.928p
Rs 1 N3 0.1
L1 N3 2 2.2u
.ends 2512_74405024022_2.2u
*******
.subckt 2512_74405024033_3.3u 1 2
Rp 1 2 2593
Cp 1 2 6.966p
Rs 1 N3 0.136
L1 N3 2 3.3u
.ends 2512_74405024033_3.3u
*******
.subckt 2512_74405024047_4.7u 1 2
Rp 1 2 3986
Cp 1 2 6.962p
Rs 1 N3 0.225
L1 N3 2 4.7u
.ends 2512_74405024047_4.7u
*******
.subckt 2512_74405024100_10u 1 2
Rp 1 2 7534
Cp 1 2 7.589p
Rs 1 N3 0.435
L1 N3 2 10u
.ends 2512_74405024100_10u
*******
.subckt 3012_744050310047_0.47u 1 2
Rp 1 2 836
Cp 1 2 3.831p
Rs 1 N3 0.028
L1 N3 2 0.47u
.ends 3012_744050310047_0.47u
*******
.subckt 3012_74405031010_1u 1 2
Rp 1 2 1251
Cp 1 2 5.888p
Rs 1 N3 0.045
L1 N3 2 1u
.ends 3012_74405031010_1u
*******
.subckt 3012_74405031015_1.5u 1 2
Rp 1 2 1524
Cp 1 2 5.275p
Rs 1 N3 0.064
L1 N3 2 1.5u
.ends 3012_74405031015_1.5u
*******
.subckt 3012_74405031022_2.2u 1 2
Rp 1 2 2126
Cp 1 2 5.715p
Rs 1 N3 0.09
L1 N3 2 2.2u
.ends 3012_74405031022_2.2u
*******
.subckt 3012_74405031033_3.3u 1 2
Rp 1 2 2811
Cp 1 2 5.52p
Rs 1 N3 0.129
L1 N3 2 3.3u
.ends 3012_74405031033_3.3u
*******
.subckt 3012_74405031047_4.7u 1 2
Rp 1 2 4435
Cp 1 2 6.438p
Rs 1 N3 0.196
L1 N3 2 4.7u
.ends 3012_74405031047_4.7u
*******
.subckt 3012_74405031100_10u 1 2
Rp 1 2 7640
Cp 1 2 5.603p
Rs 1 N3 0.395
L1 N3 2 10u
.ends 3012_74405031100_10u
*******
.subckt 4020_744050420047_0.47u 1 2
Rp 1 2 944
Cp 1 2 6.657p
Rs 1 N3 0.018
L1 N3 2 0.47u
.ends 4020_744050420047_0.47u
*******
.subckt 4020_74405042010_1u 1 2
Rp 1 2 1143
Cp 1 2 8.295p
Rs 1 N3 0.022
L1 N3 2 1u
.ends 4020_74405042010_1u
*******
.subckt 4020_74405042015_1.5u 1 2
Rp 1 2 1850
Cp 1 2 8.521p
Rs 1 N3 0.03
L1 N3 2 1.5u
.ends 4020_74405042015_1.5u
*******
.subckt 4020_74405042022_2.2u 1 2
Rp 1 2 2124
Cp 1 2 9.121p
Rs 1 N3 0.04
L1 N3 2 2.2u
.ends 4020_74405042022_2.2u
*******
.subckt 4020_74405042033_3.3u 1 2
Rp 1 2 961
Cp 1 2 39.05p
Rs 1 N3 0.06
L1 N3 2 3.3u
.ends 4020_74405042033_3.3u
*******
.subckt 4020_74405042047_4.7u 1 2
Rp 1 2 3995
Cp 1 2 9.023p
Rs 1 N3 0.09
L1 N3 2 4.7u
.ends 4020_74405042047_4.7u
*******
.subckt 4020_74405042068_6.8u 1 2
Rp 1 2 5154
Cp 1 2 10.556p
Rs 1 N3 0.13
L1 N3 2 6.8u
.ends 4020_74405042068_6.8u
*******
.subckt 4020_74405042100_10u 1 2
Rp 1 2 7441
Cp 1 2 10.21p
Rs 1 N3 0.18
L1 N3 2 10u
.ends 4020_74405042100_10u
*******
