**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  Film Capacitors
* Matchcode:              WCAP-FTXH
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/21/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 890414025007CS_33nF 1 2
Rser 1 3 0.02
Lser 2 4 8.293975014E-09
C1 3 4 0.000000033
Rpar 3 4 25000000000
.ends 890414025007CS_33nF
*******
.subckt 890414025001CS_100nF 1 2
Rser 1 3 0.0622459836403
Lser 2 4 9.907151555E-09
C1 3 4 0.0000001
Rpar 3 4 25000000000
.ends 890414025001CS_100nF
*******
.subckt 890414025008CS_120nF 1 2
Rser 1 3 0.0575
Lser 2 4 0.000000008
C1 3 4 0.00000012
Rpar 3 4 25000000000
.ends 890414025008CS_120nF
*******
.subckt 890414025002CS_150nF 1 2
Rser 1 3 0.052
Lser 2 4 0.0000000067
C1 3 4 0.00000015
Rpar 3 4 25000000000
.ends 890414025002CS_150nF
*******
.subckt 890414025003CS_220nF 1 2
Rser 1 3 0.04474
Lser 2 4 0.00000000656
C1 3 4 0.00000022
Rpar 3 4 25000000000
.ends 890414025003CS_220nF
*******
.subckt 890414025009CS_270nF 1 2
Rser 1 3 0.037
Lser 2 4 0.0000000082
C1 3 4 0.00000027
Rpar 3 4 25000000000
.ends 890414025009CS_270nF
*******
.subckt 890414025005CS_390nF 1 2
Rser 1 3 0.0315
Lser 2 4 0.000000008
C1 3 4 0.00000039
Rpar 3 4 19230000000
.ends 890414025005CS_390nF
*******
.subckt 890414025013CS_270nF 1 2
Rser 1 3 0.03083
Lser 2 4 0.00000000871
C1 3 4 0.00000027
Rpar 3 4 25000000000
.ends 890414025013CS_270nF
*******
.subckt 890414025011CS_330nF 1 2
Rser 1 3 0.03178
Lser 2 4 0.00000000834
C1 3 4 0.00000033
Rpar 3 4 25000000000
.ends 890414025011CS_330nF
*******
.subckt 890414025010CS_560nF 1 2
Rser 1 3 0.0247421343301
Lser 2 4 8.450048099E-09
C1 3 4 0.00000056
Rpar 3 4 13390000000
.ends 890414025010CS_560nF
*******
.subckt 890414025012CS_470nF 1 2
Rser 1 3 0.02693
Lser 2 4 0.00000000791
C1 3 4 0.00000047
Rpar 3 4 15950000000
.ends 890414025012CS_470nF
*******
.subckt 890414026001CS_330nF 1 2
Rser 1 3 0.046
Lser 2 4 9.360871175E-09
C1 3 4 0.00000033
Rpar 3 4 25000000000
.ends 890414026001CS_330nF
*******
.subckt 890414026002CS_390nF 1 2
Rser 1 3 0.06
Lser 2 4 0.00000001195
C1 3 4 0.00000039
Rpar 3 4 19230000000
.ends 890414026002CS_390nF
*******
.subckt 890414026003CS_470nF 1 2
Rser 1 3 0.0394787517849
Lser 2 4 9.054111549E-09
C1 3 4 0.00000047
Rpar 3 4 15950000000
.ends 890414026003CS_470nF
*******
.subckt 890414026004CS_560nF 1 2
Rser 1 3 0.0364321216625
Lser 2 4 1.1628784093E-08
C1 3 4 0.00000056
Rpar 3 4 13390000000
.ends 890414026004CS_560nF
*******
.subckt 890414026005CS_680nF 1 2
Rser 1 3 0.040848499856
Lser 2 4 1.1846559881E-08
C1 3 4 0.00000068
Rpar 3 4 11020000000
.ends 890414026005CS_680nF
*******
.subckt 890414026008CS_1.2uF 1 2
Rser 1 3 0.045
Lser 2 4 0.00000001336
C1 3 4 0.0000012
Rpar 3 4 6250000000
.ends 890414026008CS_1.2uF
*******
.subckt 890414026009CS_1.5uF 1 2
Rser 1 3 0.0258997562049
Lser 2 4 1.4071119672E-08
C1 3 4 0.0000015
Rpar 3 4 5000000000
.ends 890414026009CS_1.5uF
*******
.subckt 890414026010CS_1.8uF 1 2
Rser 1 3 0.025
Lser 2 4 0.0000000126
C1 3 4 0.0000018
Rpar 3 4 4160000000
.ends 890414026010CS_1.8uF
*******
.subckt 890414026013CS_1.2uF 1 2
Rser 1 3 0.02689
Lser 2 4 0.00000001344
C1 3 4 0.0000012
Rpar 3 4 6250000000
.ends 890414026013CS_1.2uF
*******
.subckt 890414026011CS_2.2uF 1 2
Rser 1 3 0.0236990619526
Lser 2 4 1.2406627575E-08
C1 3 4 0.0000022
Rpar 3 4 3400000000
.ends 890414026011CS_2.2uF
*******
.subckt 890414026006CS_820nF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000089
C1 3 4 0.00000082
Rpar 3 4 9140000000
.ends 890414026006CS_820nF
*******
.subckt 890414026007CS_1uF 1 2
Rser 1 3 0.0314606793523
Lser 2 4 9.186846689E-09
C1 3 4 0.000001
Rpar 3 4 7500000000
.ends 890414026007CS_1uF
*******
.subckt 890414026014CS_1uF 1 2
Rser 1 3 0.02747
Lser 2 4 0.00000001117
C1 3 4 0.000001
Rpar 3 4 7500000000
.ends 890414026014CS_1uF
*******
.subckt 890414027005CS_680nF 1 2
Rser 1 3 0.034
Lser 2 4 1.4534392213E-08
C1 3 4 0.00000068
Rpar 3 4 11020000000
.ends 890414027005CS_680nF
*******
.subckt 890414027006CS_820nF 1 2
Rser 1 3 0.0416563089983
Lser 2 4 1.3459519897E-08
C1 3 4 0.00000082
Rpar 3 4 9140000000
.ends 890414027006CS_820nF
*******
.subckt 890414027007CS_1uF 1 2
Rser 1 3 0.0396032054977
Lser 2 4 1.6648735388E-08
C1 3 4 0.000001
Rpar 3 4 7500000000
.ends 890414027007CS_1uF
*******
.subckt 890414027008CS_1.2uF 1 2
Rser 1 3 0.031
Lser 2 4 0.0000000125
C1 3 4 0.0000012
Rpar 3 4 6250000000
.ends 890414027008CS_1.2uF
*******
.subckt 890414027001CS_2.2uF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000126
C1 3 4 0.0000022
Rpar 3 4 3400000000
.ends 890414027001CS_2.2uF
*******
.subckt 890414027004CS_560nF 1 2
Rser 1 3 0.0531188513038
Lser 2 4 1.2505387039E-08
C1 3 4 0.00000056
Rpar 3 4 13390000000
.ends 890414027004CS_560nF
*******
.subckt 890414027013CS_1.2uF 1 2
Rser 1 3 0.02886
Lser 2 4 0.00000001239
C1 3 4 0.0000012
Rpar 3 4 6250000000
.ends 890414027013CS_1.2uF
*******
.subckt 890414027012CS_1uF 1 2
Rser 1 3 0.03183
Lser 2 4 0.00000001533
C1 3 4 0.000001
Rpar 3 4 7500000000
.ends 890414027012CS_1uF
*******
.subckt 890414027009CS_1.5uF 1 2
Rser 1 3 0.0308013693837
Lser 2 4 1.3622491082E-08
C1 3 4 0.0000015
Rpar 3 4 5000000000
.ends 890414027009CS_1.5uF
*******
.subckt 890414027010CS_1.8uF 1 2
Rser 1 3 0.027945366249
Lser 2 4 1.1387619177E-08
C1 3 4 0.0000018
Rpar 3 4 4160000000
.ends 890414027010CS_1.8uF
*******
.subckt 890414027014CS_1.8uF 1 2
Rser 1 3 0.02576
Lser 2 4 0.00000001407
C1 3 4 0.0000018
Rpar 3 4 4160000000
.ends 890414027014CS_1.8uF
*******
.subckt 890414027011CS_2.2uF 1 2
Rser 1 3 0.02257
Lser 2 4 0.00000001572
C1 3 4 0.0000022
Rpar 3 4 3400000000
.ends 890414027011CS_2.2uF
*******
.subckt 890414027002CS_3.3uF 1 2
Rser 1 3 0.0222982936209
Lser 2 4 1.3650736089E-08
C1 3 4 0.0000033
Rpar 3 4 2270000000
.ends 890414027002CS_3.3uF
*******
.subckt 890414027003CS_4.7uF 1 2
Rser 1 3 0.020284320757
Lser 2 4 1.2805463076E-08
C1 3 4 0.0000047
Rpar 3 4 1590000000
.ends 890414027003CS_4.7uF
*******
.subckt 890414028005CS_3.3uF 1 2
Rser 1 3 0.02191
Lser 2 4 0.00000001686
C1 3 4 0.0000033
Rpar 3 4 2270000000
.ends 890414028005CS_3.3uF
*******
.subckt 890414028001CS_4.7uF 1 2
Rser 1 3 0.0181533724788
Lser 2 4 1.8406086695E-08
C1 3 4 0.0000047
Rpar 3 4 1590000000
.ends 890414028001CS_4.7uF
*******
.subckt 890414028006CS_4.7uF 1 2
Rser 1 3 0.01576
Lser 2 4 0.00000001962
C1 3 4 0.0000047
Rpar 3 4 1590000000
.ends 890414028006CS_4.7uF
*******
.subckt 890414028003CS_6.8uF 1 2
Rser 1 3 0.0152571553588
Lser 2 4 1.6120022101E-08
C1 3 4 0.0000068
Rpar 3 4 1100000000
.ends 890414028003CS_6.8uF
*******
.subckt 890414028002CS_10uF 1 2
Rser 1 3 0.0112884501567
Lser 2 4 2.3263893093E-08
C1 3 4 0.00001
Rpar 3 4 750000000
.ends 890414028002CS_10uF
*******
.subckt 890414028007CS_10uF 1 2
Rser 1 3 0.01079
Lser 2 4 0.00000002214
C1 3 4 0.00001
Rpar 3 4 750000000
.ends 890414028007CS_10uF
*******
