**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT High Current Cube Inductor
* Matchcode:             WE-HCC
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/9/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1090_7443330022_0.22u 1 2
Rp 1 2 332.13
Cp 1 2 1.27930787427177p
Rs 1 N3 0.0014
L1 N3 2 0.22u
.ends 1090_7443330022_0.22u
*******
.subckt 1090_7443330033_0.33u 1 2
Rp 1 2 324.68
Cp 1 2 1.27327909069839p
Rs 1 N3 0.0014
L1 N3 2 0.3183u
.ends 1090_7443330033_0.33u
*******
.subckt 1090_7443330047_0.47u 1 2
Rp 1 2 532.74
Cp 1 2 1.93708826156436p
Rs 1 N3 0.0016
L1 N3 2 0.5108u
.ends 1090_7443330047_0.47u
*******
.subckt 1090_7443330068_0.68u 1 2
Rp 1 2 834.55
Cp 1 2 1.77259290647684p
Rs 1 N3 0.00215
L1 N3 2 0.72908u
.ends 1090_7443330068_0.68u
*******
.subckt 1090_7443330082_0.82u 1 2
Rp 1 2 824.42
Cp 1 2 2.2135025319605p
Rs 1 N3 0.00215
L1 N3 2 0.79469u
.ends 1090_7443330082_0.82u
*******
.subckt 1090_7443330100_1u 1 2
Rp 1 2 803.92
Cp 1 2 2.061p
Rs 1 N3 0.00215
L1 N3 2 1.123u
.ends 1090_7443330100_1u
*******
.subckt 1090_7443330150_1.5u 1 2
Rp 1 2 1327
Cp 1 2 2.64p
Rs 1 N3 0.00335
L1 N3 2 1.533u
.ends 1090_7443330150_1.5u
*******
.subckt 1090_7443330220_2.2u 1 2
Rp 1 2 1784
Cp 1 2 1.727p
Rs 1 N3 0.0046
L1 N3 2 1.945u
.ends 1090_7443330220_2.2u
*******
.subckt 1090_7443330330_3.3u 1 2
Rp 1 2 2701
Cp 1 2 2.959p
Rs 1 N3 0.0065
L1 N3 2 3.243u
.ends 1090_7443330330_3.3u
*******
.subckt 1090_7443330470_4.7u 1 2
Rp 1 2 3350
Cp 1 2 2.442p
Rs 1 N3 0.0094
L1 N3 2 4.216u
.ends 1090_7443330470_4.7u
*******
.subckt 1090_7443330680_6.8u 1 2
Rp 1 2 4635
Cp 1 2 2.114p
Rs 1 N3 0.01415
L1 N3 2 6.255u
.ends 1090_7443330680_6.8u
*******
.subckt 1090_7443330820_8.2u 1 2
Rp 1 2 4441.2
Cp 1 2 2.933p
Rs 1 N3 0.01415
L1 N3 2 8.195u
.ends 1090_7443330820_8.2u
*******
.subckt 1090_7443331000_10u 1 2
Rp 1 2 5570
Cp 1 2 2.139p
Rs 1 N3 0.02275
L1 N3 2 9.378u
.ends 1090_7443331000_10u
*******
.subckt 1210_7443320022_0.22u 1 2
Rp 1 2 292.2
Cp 1 2 1.81044846783251p
Rs 1 N3 0.0011
L1 N3 2 0.20697u
.ends 1210_7443320022_0.22u
*******
.subckt 1210_7443310022_0.22u 1 2
Rp 1 2 158.8
Cp 1 2 2.87844271711149p
Rs 1 N3 0.0011
L1 N3 2 0.22u
.ends 1210_7443310022_0.22u
*******
.subckt 1210_7443320033_0.33u 1 2
Rp 1 2 305.62
Cp 1 2 1.83824609644555p
Rs 1 N3 0.0011
L1 N3 2 0.34449u
.ends 1210_7443320033_0.33u
*******
.subckt 1210_7443310033_0.33u 1 2
Rp 1 2 136.36
Cp 1 2 2.36908865605884p
Rs 1 N3 0.0011
L1 N3 2 0.33u
.ends 1210_7443310033_0.33u
*******
.subckt 1210_7443320047_0.47u 1 2
Rp 1 2 546.64
Cp 1 2 2.47154979003109p
Rs 1 N3 0.00135
L1 N3 2 0.4555u
.ends 1210_7443320047_0.47u
*******
.subckt 1210_7443310047_0.47u 1 2
Rp 1 2 166.88
Cp 1 2 5.38942466182577p
Rs 1 N3 0.00135
L1 N3 2 0.47u
.ends 1210_7443310047_0.47u
*******
.subckt 1210_7443320068_0.68u 1 2
Rp 1 2 514.54
Cp 1 2 2.87083500434996p
Rs 1 N3 0.00135
L1 N3 2 0.7292u
.ends 1210_7443320068_0.68u
*******
.subckt 1210_7443310068_0.68u 1 2
Rp 1 2 135.24
Cp 1 2 2.58683577518189p
Rs 1 N3 0.00135
L1 N3 2 0.68u
.ends 1210_7443310068_0.68u
*******
.subckt 1210_7443320082_0.82u 1 2
Rp 1 2 783.38
Cp 1 2 2.82294616188355p
Rs 1 N3 0.00185
L1 N3 2 0.8973u
.ends 1210_7443320082_0.82u
*******
.subckt 1210_7443310082_0.82u 1 2
Rp 1 2 253.76
Cp 1 2 3.42278169185611p
Rs 1 N3 0.00195
L1 N3 2 0.82u
.ends 1210_7443310082_0.82u
*******
.subckt 1210_7443320100_1u 1 2
Rp 1 2 782.48
Cp 1 2 2.66794770657985p
Rs 1 N3 0.00185
L1 N3 2 1.052u
.ends 1210_7443320100_1u
*******
.subckt 1210_7443310100_1u 1 2
Rp 1 2 146.9
Cp 1 2 2.09341288517199p
Rs 1 N3 0.00195
L1 N3 2 1u
.ends 1210_7443310100_1u
*******
.subckt 1210_7443320150_1.5u 1 2
Rp 1 2 1232
Cp 1 2 2.426244504791p
Rs 1 N3 0.00295
L1 N3 2 1.445u
.ends 1210_7443320150_1.5u
*******
.subckt 1210_7443310150_1.5u 1 2
Rp 1 2 176.09
Cp 1 2 2.08479801733178p
Rs 1 N3 0.0028
L1 N3 2 1.5u
.ends 1210_7443310150_1.5u
*******
.subckt 1210_7443320220_2.2u 1 2
Rp 1 2 1858
Cp 1 2 2.39334782842184p
Rs 1 N3 0.0039
L1 N3 2 2.505u
.ends 1210_7443320220_2.2u
*******
.subckt 1210_7443310220_2.2u 1 2
Rp 1 2 365.45
Cp 1 2 3.19826968567943p
Rs 1 N3 0.00375
L1 N3 2 2.2u
.ends 1210_7443310220_2.2u
*******
.subckt 1210_7443320330_3.3u 1 2
Rp 1 2 2269
Cp 1 2 4.74421185019874p
Rs 1 N3 0.0052
L1 N3 2 3.337u
.ends 1210_7443320330_3.3u
*******
.subckt 1210_7443310330_3.3u 1 2
Rp 1 2 344.22
Cp 1 2 12.281355593009p
Rs 1 N3 0.00695
L1 N3 2 3.3u
.ends 1210_7443310330_3.3u
*******
.subckt 1210_7443310390_3.9u 1 2
Rp 1 2 799.7
Cp 1 2 3.20738156512581p
Rs 1 N3 0.01
L1 N3 2 3.9u
.ends 1210_7443310390_3.9u
*******
.subckt 1210_7443320470_4.7u 1 2
Rp 1 2 2952
Cp 1 2 3.43787946669125p
Rs 1 N3 0.00725
L1 N3 2 4.605u
.ends 1210_7443320470_4.7u
*******
.subckt 1210_7443310470_4.7u 1 2
Rp 1 2 639.9
Cp 1 2 3.3683904136411p
Rs 1 N3 0.01
L1 N3 2 4.7u
.ends 1210_7443310470_4.7u
*******
.subckt 1210_7443320680_6.8u 1 2
Rp 1 2 2684
Cp 1 2 3.15884396273544p
Rs 1 N3 0.01015
L1 N3 2 6.546u
.ends 1210_7443320680_6.8u
*******
.subckt 1210_7443320820_8.2u 1 2
Rp 1 2 4179
Cp 1 2 2.46181781794726p
Rs 1 N3 0.0106
L1 N3 2 8.3994u
.ends 1210_7443320820_8.2u
*******
.subckt 1210_7443321000_10u 1 2
Rp 1 2 5020
Cp 1 2 4.2085642219034p
Rs 1 N3 0.01535
L1 N3 2 9.63u
.ends 1210_7443321000_10u
*******
.subckt 8070_7443340030_0.3u 1 2
Rp 1 2 470.91
Cp 1 2 1.31705685223352p
Rs 1 N3 0.0023
L1 N3 2 0.30772u
.ends 8070_7443340030_0.3u
*******
.subckt 8070_7443340047_0.47u 1 2
Rp 1 2 621.28
Cp 1 2 1.05835048459105p
Rs 1 N3 0.00265
L1 N3 2 0.38294u
.ends 8070_7443340047_0.47u
*******
.subckt 8070_7443340068_0.68u 1 2
Rp 1 2 699.24
Cp 1 2 1.32877703531752p
Rs 1 N3 0.00265
L1 N3 2 0.58836u
.ends 8070_7443340068_0.68u
*******
.subckt 8070_7443340100_1u 1 2
Rp 1 2 1166
Cp 1 2 1.31147015643337p
Rs 1 N3 0.0036
L1 N3 2 0.98543u
.ends 8070_7443340100_1u
*******
.subckt 8070_7443340150_1.5u 1 2
Rp 1 2 1584
Cp 1 2 1.389p
Rs 1 N3 0.0053
L1 N3 2 1.295u
.ends 8070_7443340150_1.5u
*******
.subckt 8070_7443340220_2.2u 1 2
Rp 1 2 1468
Cp 1 2 1.471p
Rs 1 N3 0.0053
L1 N3 2 1.97u
.ends 8070_7443340220_2.2u
*******
.subckt 8070_7443340330_3.3u 1 2
Rp 1 2 2132
Cp 1 2 1.438p
Rs 1 N3 0.0075
L1 N3 2 2.919u
.ends 8070_7443340330_3.3u
*******
.subckt 8070_7443340470_4.7u 1 2
Rp 1 2 2026
Cp 1 2 2.718p
Rs 1 N3 0.0127
L1 N3 2 4.386u
.ends 8070_7443340470_4.7u
*******
.subckt 8070_7443340680_6.8u 1 2
Rp 1 2 2891
Cp 1 2 2.779p
Rs 1 N3 0.0233
L1 N3 2 6.407u
.ends 8070_7443340680_6.8u
*******
.subckt 8070_7443341000_10u 1 2
Rp 1 2 6278
Cp 1 2 3.371p
Rs 1 N3 0.0385
L1 N3 2 8.837u
.ends 8070_7443341000_10u
*******
