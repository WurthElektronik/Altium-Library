**************************************************
* Manufacturer:          Würth Elektronik 
* Kinds:                 Multilayer Ceramic Chip Capacitors
* Matchcode:             WCAP-CSRF
* Library Type:          LTspice
* Version:               rev23a
* Created/modified by:   Ella
* Date and Time:         9/19/2023
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2023 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 0201_885392004001_0.2pF 1 2
Rser 1 3 0.5187
Lser 2 4 0.00000000058
C1 3 4 0.0000000000002
Rpar 3 4 10000000000
.ends 0201_885392004001_0.2pF
*******
.subckt 0201_885392004002_1pF 1 2
Rser 1 3 1.0325
Lser 2 4 0.000000000343
C1 3 4 0.000000000001
Rpar 3 4 10000000000
.ends 0201_885392004002_1pF
*******
.subckt 0201_885392004003_1.2pF 1 2
Rser 1 3 0.9171
Lser 2 4 0.000000000335
C1 3 4 0.0000000000012
Rpar 3 4 10000000000
.ends 0201_885392004003_1.2pF
*******
.subckt 0201_885392004004_1.5pF 1 2
Rser 1 3 0.6731
Lser 2 4 0.000000000302
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0201_885392004004_1.5pF
*******
.subckt 0201_885392004005_2.2pF 1 2
Rser 1 3 0.3893
Lser 2 4 0.000000000271
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0201_885392004005_2.2pF
*******
.subckt 0201_885392004006_2.7pF 1 2
Rser 1 3 0.3777
Lser 2 4 0.000000000352
C1 3 4 0.0000000000027
Rpar 3 4 10000000000
.ends 0201_885392004006_2.7pF
*******
.subckt 0201_885392004007_3.3pF 1 2
Rser 1 3 0.3218
Lser 2 4 0.000000000268
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0201_885392004007_3.3pF
*******
.subckt 0201_885392004008_4.7pF 1 2
Rser 1 3 0.2363
Lser 2 4 0.000000000248
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0201_885392004008_4.7pF
*******
.subckt 0201_885392004009_5.6pF 1 2
Rser 1 3 0.4286
Lser 2 4 0.000000000266
C1 3 4 0.0000000000056
Rpar 3 4 10000000000
.ends 0201_885392004009_5.6pF
*******
.subckt 0201_885392004010_9pF 1 2
Rser 1 3 0.1717
Lser 2 4 0.000000000228
C1 3 4 0.000000000009
Rpar 3 4 10000000000
.ends 0201_885392004010_9pF
*******
.subckt 0201_885392004011_33pF 1 2
Rser 1 3 0.1789
Lser 2 4 0.000000000265
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0201_885392004011_33pF
*******
.subckt 0402_885392005001_0.3pF 1 2
Rser 1 3 0.61864
Lser 2 4 0.00000000063
C1 3 4 0.0000000000003
Rpar 3 4 10000000000
.ends 0402_885392005001_0.3pF
*******
.subckt 0402_885392005002_0.4pF 1 2
Rser 1 3 0.818
Lser 2 4 0.000000000314
C1 3 4 0.0000000000004
Rpar 3 4 10000000000
.ends 0402_885392005002_0.4pF
*******
.subckt 0402_885392005003_0.4pF 1 2
Rser 1 3 1.186
Lser 2 4 0.000000000342
C1 3 4 0.0000000000004
Rpar 3 4 10000000000
.ends 0402_885392005003_0.4pF
*******
.subckt 0402_885392005004_0.5pF 1 2
Rser 1 3 0.7967
Lser 2 4 0.000000000378
C1 3 4 0.0000000000005
Rpar 3 4 10000000000
.ends 0402_885392005004_0.5pF
*******
.subckt 0402_885392005005_1pF 1 2
Rser 1 3 1.1161
Lser 2 4 0.000000000448
C1 3 4 0.000000000001
Rpar 3 4 10000000000
.ends 0402_885392005005_1pF
*******
.subckt 0402_885392005006_1pF 1 2
Rser 1 3 1.2856
Lser 2 4 0.000000000401
C1 3 4 0.000000000001
Rpar 3 4 10000000000
.ends 0402_885392005006_1pF
*******
.subckt 0402_885392005007_1.5pF 1 2
Rser 1 3 1.001
Lser 2 4 0.000000000414
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0402_885392005007_1.5pF
*******
.subckt 0402_885392005008_1.8pF 1 2
Rser 1 3 0.4527
Lser 2 4 0.000000000392
C1 3 4 0.0000000000018
Rpar 3 4 10000000000
.ends 0402_885392005008_1.8pF
*******
.subckt 0402_885392005009_2.3pF 1 2
Rser 1 3 0.8313
Lser 2 4 0.000000000332
C1 3 4 0.0000000000023
Rpar 3 4 10000000000
.ends 0402_885392005009_2.3pF
*******
.subckt 0402_885392005010_3pF 1 2
Rser 1 3 0.771
Lser 2 4 0.000000000307
C1 3 4 0.000000000003
Rpar 3 4 10000000000
.ends 0402_885392005010_3pF
*******
.subckt 0402_885392005011_3.3pF 1 2
Rser 1 3 0.5129
Lser 2 4 0.000000000385
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0402_885392005011_3.3pF
*******
.subckt 0402_885392005012_4.7pF 1 2
Rser 1 3 0.4028
Lser 2 4 0.000000000404
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0402_885392005012_4.7pF
*******
.subckt 0402_885392005013_5.6pF 1 2
Rser 1 3 0.6213
Lser 2 4 0.000000000335
C1 3 4 0.0000000000056
Rpar 3 4 10000000000
.ends 0402_885392005013_5.6pF
*******
.subckt 0402_885392005014_9pF 1 2
Rser 1 3 0.2845
Lser 2 4 0.000000000364
C1 3 4 0.000000000009
Rpar 3 4 10000000000
.ends 0402_885392005014_9pF
*******
.subckt 0402_885392005019_0.7pF 1 2
Rser 1 3 1.3365
Lser 2 4 0.000000000388
C1 3 4 0.0000000000007
Rpar 3 4 10000000000
.ends 0402_885392005019_0.7pF
*******
.subckt 0402_885392005022_0.9pF 1 2
Rser 1 3 0.7061
Lser 2 4 0.00000000036
C1 3 4 0.0000000000009
Rpar 3 4 10000000000
.ends 0402_885392005022_0.9pF
*******
.subckt 0402_885392005024_1.2pF 1 2
Rser 1 3 0.4162
Lser 2 4 0.000000000378
C1 3 4 0.0000000000012
Rpar 3 4 10000000000
.ends 0402_885392005024_1.2pF
*******
.subckt 0402_885392005030_2pF 1 2
Rser 1 3 1.049
Lser 2 4 0.000000000287
C1 3 4 0.000000000002
Rpar 3 4 10000000000
.ends 0402_885392005030_2pF
*******
.subckt 0402_885392005032_2.2pF 1 2
Rser 1 3 1.0061
Lser 2 4 0.000000000362
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0402_885392005032_2.2pF
*******
.subckt 0402_885392005034_2.4pF 1 2
Rser 1 3 0.4264
Lser 2 4 0.000000000298
C1 3 4 0.0000000000024
Rpar 3 4 10000000000
.ends 0402_885392005034_2.4pF
*******
.subckt 0402_885392005037_2.7pF 1 2
Rser 1 3 0.315
Lser 2 4 0.000000000276
C1 3 4 0.0000000000027
Rpar 3 4 10000000000
.ends 0402_885392005037_2.7pF
*******
.subckt 0402_885392005044_3.6pF 1 2
Rser 1 3 0.249
Lser 2 4 0.00000000027
C1 3 4 0.0000000000036
Rpar 3 4 10000000000
.ends 0402_885392005044_3.6pF
*******
.subckt 0402_885392005047_3.9pF 1 2
Rser 1 3 0.5269
Lser 2 4 0.000000000286
C1 3 4 0.0000000000039
Rpar 3 4 10000000000
.ends 0402_885392005047_3.9pF
*******
.subckt 0402_885392005051_4.3pF 1 2
Rser 1 3 0.853
Lser 2 4 0.000000000407
C1 3 4 0.0000000000043
Rpar 3 4 10000000000
.ends 0402_885392005051_4.3pF
*******
.subckt 0402_885392005074_6.8pF 1 2
Rser 1 3 0.3481
Lser 2 4 0.000000000353
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0402_885392005074_6.8pF
*******
.subckt 0402_885392005081_7.5pF 1 2
Rser 1 3 0.2387
Lser 2 4 0.000000000381
C1 3 4 0.0000000000075
Rpar 3 4 10000000000
.ends 0402_885392005081_7.5pF
*******
.subckt 0402_885392005088_8.2pF 1 2
Rser 1 3 0.3077
Lser 2 4 0.000000000518
C1 3 4 0.0000000000082
Rpar 3 4 10000000000
.ends 0402_885392005088_8.2pF
*******
.subckt 0402_885392005097_9.1pF 1 2
Rser 1 3 0.7892
Lser 2 4 0.000000000379
C1 3 4 0.0000000000091
Rpar 3 4 10000000000
.ends 0402_885392005097_9.1pF
*******
.subckt 0402_885392005106_10pF 1 2
Rser 1 3 0.493
Lser 2 4 0.000000000305
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885392005106_10pF
*******
.subckt 0402_885392005110_15pF 1 2
Rser 1 3 0.2685
Lser 2 4 0.000000000398
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885392005110_15pF
*******
.subckt 0402_885392005114_22pF 1 2
Rser 1 3 0.2703
Lser 2 4 0.000000000328
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885392005114_22pF
*******
.subckt 0402_885392005116_27pF 1 2
Rser 1 3 0.2206
Lser 2 4 0.000000000478
C1 3 4 0.000000000027
Rpar 3 4 10000000000
.ends 0402_885392005116_27pF
*******
.subckt 0402_885392005127_12pF 1 2
Rser 1 3 0.4176
Lser 2 4 0.00000000033
C1 3 4 0.000000000012
Rpar 3 4 10000000000
.ends 0402_885392005127_12pF
*******
.subckt 0402_885392005130_0.8pF 1 2
Rser 1 3 0.3869
Lser 2 4 0.000000000328
C1 3 4 0.0000000000008
Rpar 3 4 10000000000
.ends 0402_885392005130_0.8pF
*******
