**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ASLU
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         5/31/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 865090140001_10uF 1 2
Rser 1 3 2.31804872278
Lser 2 4 1.92353053E-09
C1 3 4 0.00001
Rpar 3 4 2100000
.ends 865090140001_10uF
*******
.subckt 865090140002_22uF 1 2
Rser 1 3 2.43004421152
Lser 2 4 1.073688846E-09
C1 3 4 0.000022
Rpar 3 4 2100000
.ends 865090140002_22uF
*******
.subckt 865090140003_33uF 1 2
Rser 1 3 2.03800634474
Lser 2 4 1.926725732E-09
C1 3 4 0.000033
Rpar 3 4 2100000
.ends 865090140003_33uF
*******
.subckt 865090140004_47uF 1 2
Rser 1 3 2.40992855164
Lser 2 4 1.851137929E-09
C1 3 4 0.000047
Rpar 3 4 2100000
.ends 865090140004_47uF
*******
.subckt 865090142005_100uF 1 2
Rser 1 3 0.59
Lser 2 4 0.00000000002
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865090142005_100uF
*******
.subckt 865090145006_220uF 1 2
Rser 1 3 0.53259101206
Lser 2 4 4.360458939E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545454
.ends 865090145006_220uF
*******
.subckt 865090145008_330uF 1 2
Rser 1 3 0.3
Lser 2 4 0.00000000008
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865090145008_330uF
*******
.subckt 865090149007_220uF 1 2
Rser 1 3 0.34
Lser 2 4 0.00000000012
C1 3 4 0.00022
Rpar 3 4 454545.454545454
.ends 865090149007_220uF
*******
.subckt 865090149009_330uF 1 2
Rser 1 3 0.361
Lser 2 4 3.67826263073994E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865090149009_330uF
*******
.subckt 865090168010_22uF 1 2
Rser 1 3 1.95
Lser 2 4 0.00000000000007
C1 3 4 0.000022
Rpar 3 4 2100000
.ends 865090168010_22uF
*******
.subckt 865090240001_10uF 1 2
Rser 1 3 2.46985323746
Lser 2 4 9.42355697E-10
C1 3 4 0.00001
Rpar 3 4 3333333.33333333
.ends 865090240001_10uF
*******
.subckt 865090240002_22uF 1 2
Rser 1 3 2.59906374467
Lser 2 4 8.19894981E-10
C1 3 4 0.000022
Rpar 3 4 3333333.33333333
.ends 865090240002_22uF
*******
.subckt 865090242003_33uF 1 2
Rser 1 3 1.54226230476
Lser 2 4 2.423178826E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865090242003_33uF
*******
.subckt 865090243004_47uF 1 2
Rser 1 3 0.976158717401
Lser 2 4 3.326744982E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865090243004_47uF
*******
.subckt 865090245005_100uF 1 2
Rser 1 3 0.481799881175
Lser 2 4 4.286638938E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865090245005_100uF
*******
.subckt 865090245007_220uF 1 2
Rser 1 3 0.5
Lser 2 4 0.00000000014
C1 3 4 0.000047
Rpar 3 4 454545.454545455
.ends 865090245007_220uF
*******
.subckt 865090249006_100uF 1 2
Rser 1 3 0.662722204299
Lser 2 4 3.76317886E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865090249006_100uF
*******
.subckt 865090249008_220uF 1 2
Rser 1 3 0.571673841911
Lser 2 4 5.782497809E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865090249008_220uF
*******
.subckt 865090268009_10uF 1 2
Rser 1 3 2.05
Lser 2 4 0.00000000000023
C1 3 4 0.00001
Rpar 3 4 3333333.33333333
.ends 865090268009_10uF
*******
.subckt 865090340001_4.7uF 1 2
Rser 1 3 2.00437098761
Lser 2 4 8.90117854E-10
C1 3 4 0.0000047
Rpar 3 4 5333333.33333333
.ends 865090340001_4.7uF
*******
.subckt 865090340002_10uF 1 2
Rser 1 3 1.45
Lser 2 4 0.0000000000013
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 865090340002_10uF
*******
.subckt 865090342003_22uF 1 2
Rser 1 3 1.2
Lser 2 4 1.742530489E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865090342003_22uF
*******
.subckt 865090343004_33uF 1 2
Rser 1 3 0.65
Lser 2 4 0.000000002245
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865090343004_33uF
*******
.subckt 865090343005_47uF 1 2
Rser 1 3 0.98
Lser 2 4 0.000000002427
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865090343005_47uF
*******
.subckt 865090345006_100uF 1 2
Rser 1 3 0.36
Lser 2 4 0.000000002663
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865090345006_100uF
*******
.subckt 865090349007_100uF 1 2
Rser 1 3 0.362
Lser 2 4 2.07208082969975E-08
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865090349007_100uF
*******
.subckt 865090368008_10uF 1 2
Rser 1 3 2
Lser 2 4 0.00000000000018
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 865090368008_10uF
*******
.subckt 865090440001_3.3uF 1 2
Rser 1 3 2.49490253618
Lser 2 4 1.57762562E-09
C1 3 4 0.0000033
Rpar 3 4 8333333.33333333
.ends 865090440001_3.3uF
*******
.subckt 865090440002_4.7uF 1 2
Rser 1 3 1.92921464604
Lser 2 4 0.0000000005517
C1 3 4 0.0000047
Rpar 3 4 8333333.33333333
.ends 865090440002_4.7uF
*******
.subckt 865090440003_10uF 1 2
Rser 1 3 2.22516828923
Lser 2 4 0.00000000083491
C1 3 4 0.00001
Rpar 3 4 8333333.33333333
.ends 865090440003_10uF
*******
.subckt 865090442004_22uF 1 2
Rser 1 3 1.87747357625
Lser 2 4 1.038862593E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865090442004_22uF
*******
.subckt 865090443005_33uF 1 2
Rser 1 3 1.15439703162
Lser 2 4 2.38622471E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865090443005_33uF
*******
.subckt 865090445006_47uF 1 2
Rser 1 3 0.68986
Lser 2 4 2.85216443E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865090445006_47uF
*******
.subckt 865090445008_100uF 1 2
Rser 1 3 0.5
Lser 2 4 0.0000000029
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865090445008_100uF
*******
.subckt 865090449007_47uF 1 2
Rser 1 3 0.5
Lser 2 4 0.00000000014
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865090449007_47uF
*******
.subckt 865090449009_100uF 1 2
Rser 1 3 0.55427
Lser 2 4 3.868433908E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865090449009_100uF
*******
.subckt 865090468010_3.3uF 1 2
Rser 1 3 2.1
Lser 2 4 0.00000000000045
C1 3 4 0.0000033
Rpar 3 4 8333333.33333333
.ends 865090468010_3.3uF
*******
.subckt 865090468011_4.7uF 1 2
Rser 1 3 2.2
Lser 2 4 0.0000000000002
C1 3 4 0.0000047
Rpar 3 4 8333333.33333333
.ends 865090468011_4.7uF
*******
.subckt 865090540002_3.3uF 1 2
Rser 1 3 2.57363294267
Lser 2 4 1.847982175E-09
C1 3 4 0.0000033
Rpar 3 4 11666666.6666667
.ends 865090540002_3.3uF
*******
.subckt 865090543004_10uF 1 2
Rser 1 3 0.923049824619
Lser 2 4 3.698328149E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865090543004_10uF
*******
.subckt 865090543005_22uF 1 2
Rser 1 3 1.64444076348
Lser 2 4 3.600545602E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 865090543005_22uF
*******
.subckt 865090545006_33uF 1 2
Rser 1 3 0.715670650228
Lser 2 4 4.7196452E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865090545006_33uF
*******
.subckt 865090545008_47uF 1 2
Rser 1 3 0.757598567578
Lser 2 4 4.004967921E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865090545008_47uF
*******
.subckt 865090549007_33uF 1 2
Rser 1 3 0.55
Lser 2 4 0.00000000022
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865090549007_33uF
*******
.subckt 865090549009_47uF 1 2
Rser 1 3 0.779962845375
Lser 2 4 5.951668821E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865090549009_47uF
*******
.subckt 865090640001_100nF 1 2
Rser 1 3 1.44131674907
Lser 2 4 2.465045867E-09
C1 3 4 0.0000001
Rpar 3 4 16666666.6666667
.ends 865090640001_100nF
*******
.subckt 865090640002_220nF 1 2
Rser 1 3 1.8778458778
Lser 2 4 2.008178176E-09
C1 3 4 0.00000022
Rpar 3 4 16666666.6666667
.ends 865090640002_220nF
*******
.subckt 865090640003_330nF 1 2
Rser 1 3 1.8433070224
Lser 2 4 2.23671331E-09
C1 3 4 0.00000033
Rpar 3 4 16666666.6666667
.ends 865090640003_330nF
*******
.subckt 865090640004_470nF 1 2
Rser 1 3 1.68358622089
Lser 2 4 2.187302537E-09
C1 3 4 0.00000047
Rpar 3 4 16666666.6666667
.ends 865090640004_470nF
*******
.subckt 865090640005_1uF 1 2
Rser 1 3 1.5
Lser 2 4 0.0000000000014
C1 3 4 0.000001
Rpar 3 4 16666666.6666667
.ends 865090640005_1uF
*******
.subckt 865090640006_2.2uF 1 2
Rser 1 3 2.19211655403
Lser 2 4 1.369422771E-09
C1 3 4 0.0000022
Rpar 3 4 16666666.6666667
.ends 865090640006_2.2uF
*******
.subckt 865090640007_3.3uF 1 2
Rser 1 3 2.51273779765
Lser 2 4 1.835347864E-09
C1 3 4 0.0000033
Rpar 3 4 16666666.6666667
.ends 865090640007_3.3uF
*******
.subckt 865090643008_4.7uF 1 2
Rser 1 3 1.44201944388
Lser 2 4 2.242711315E-09
C1 3 4 0.0000047
Rpar 3 4 16666666.6666667
.ends 865090643008_4.7uF
*******
.subckt 865090643009_10uF 1 2
Rser 1 3 1.69799368738
Lser 2 4 2.84000955E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865090643009_10uF
*******
.subckt 865090645010_22uF 1 2
Rser 1 3 0.760152002813
Lser 2 4 3.998511065E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865090645010_22uF
*******
.subckt 865090645012_33uF 1 2
Rser 1 3 0.721220480805
Lser 2 4 4.297851511E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865090645012_33uF
*******
.subckt 865090649011_22uF 1 2
Rser 1 3 0.515
Lser 2 4 0.0000000002
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865090649011_22uF
*******
.subckt 865090649013_33uF 1 2
Rser 1 3 0.721206333687
Lser 2 4 6.186671729E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865090649013_33uF
*******
.subckt 865090668014_100nF 1 2
Rser 1 3 1.9
Lser 2 4 0.0000000000025
C1 3 4 0.0000001
Rpar 3 4 16666666.6666667
.ends 865090668014_100nF
*******
.subckt 865090668015_220nF 1 2
Rser 1 3 1.9
Lser 2 4 0.000000000002
C1 3 4 0.00000022
Rpar 3 4 16666666.6666667
.ends 865090668015_220nF
*******
.subckt 865090668016_330nF 1 2
Rser 1 3 1.9
Lser 2 4 0.0000000000007
C1 3 4 0.00000033
Rpar 3 4 16666666.6666667
.ends 865090668016_330nF
*******
.subckt 865090749001_22uF 1 2
Rser 1 3 0.43
Lser 2 4 0.0000000003
C1 3 4 0.000022
Rpar 3 4 4500000
.ends 865090749001_22uF
*******
.subckt 865090768002_100nF 1 2
Rser 1 3 1.9
Lser 2 4 0.0000000000028
C1 3 4 0.0000001
Rpar 3 4 21000000
.ends 865090768002_100nF
*******
.subckt 865090768003_220nF 1 2
Rser 1 3 2.2
Lser 2 4 1.211321E-12
C1 3 4 0.00000022
Rpar 3 4 21000000
.ends 865090768003_220nF
*******
.subckt 865090768004_330nF 1 2
Rser 1 3 1.9
Lser 2 4 0.0000000000007
C1 3 4 0.00000033
Rpar 3 4 21000000
.ends 865090768004_330nF
*******
.subckt 865090768005_470nF 1 2
Rser 1 3 2.2
Lser 2 4 0.0000000000007
C1 3 4 0.00000047
Rpar 3 4 21000000
.ends 865090768005_470nF
*******
