**************************************************
* Manufacturer:          Würth Elektronik 
* Kinds:                 Film Capacitors
* Matchcode:             WCAP-FTXX
* Library Type:          LTspice
* Version:               rev23a
* Created/modified by:   Ella
* Date and Time:         11/1/2023
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2023 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 890334022007_15nF 1 2
Rser 1 3 0.062
Lser 2 4 0.0000000039
C1 3 4 0.000000015
Rpar 3 4 30000000000
.ends 890334022007_15nF
*******
.subckt 890334022007CS_15nF 1 2
Rser 1 3 0.062
Lser 2 4 0.0000000039
C1 3 4 0.000000015
Rpar 3 4 30000000000
.ends 890334022007CS_15nF
*******
.subckt 890334022017_68nF 1 2
Rser 1 3 0.056
Lser 2 4 0.000000006
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890334022017_68nF
*******
.subckt 890334022017CS_68nF 1 2
Rser 1 3 0.056
Lser 2 4 0.000000006
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890334022017CS_68nF
*******
.subckt 890334023002_5.6nF 1 2
Rser 1 3 0.13
Lser 2 4 0.0000000057
C1 3 4 0.0000000056
Rpar 3 4 30000000000
.ends 890334023002_5.6nF
*******
.subckt 890334023002CS_5.6nF 1 2
Rser 1 3 0.13
Lser 2 4 0.0000000057
C1 3 4 0.0000000056
Rpar 3 4 30000000000
.ends 890334023002CS_5.6nF
*******
.subckt 890334023003_6.8nF 1 2
Rser 1 3 0.153
Lser 2 4 0.0000000063
C1 3 4 0.0000000068
Rpar 3 4 30000000000
.ends 890334023003_6.8nF
*******
.subckt 890334023003CS_6.8nF 1 2
Rser 1 3 0.153
Lser 2 4 0.0000000063
C1 3 4 0.0000000068
Rpar 3 4 30000000000
.ends 890334023003CS_6.8nF
*******
.subckt 890334023004_8.2nF 1 2
Rser 1 3 0.128
Lser 2 4 0.0000000061
C1 3 4 0.0000000082
Rpar 3 4 30000000000
.ends 890334023004_8.2nF
*******
.subckt 890334023004CS_8.2nF 1 2
Rser 1 3 0.128
Lser 2 4 0.0000000061
C1 3 4 0.0000000082
Rpar 3 4 30000000000
.ends 890334023004CS_8.2nF
*******
.subckt 890334023006_10nF 1 2
Rser 1 3 0.113
Lser 2 4 0.0000000072
C1 3 4 0.00000001
Rpar 3 4 30000000000
.ends 890334023006_10nF
*******
.subckt 890334023006CS_10nF 1 2
Rser 1 3 0.113
Lser 2 4 0.0000000072
C1 3 4 0.00000001
Rpar 3 4 30000000000
.ends 890334023006CS_10nF
*******
.subckt 890334023007_12nF 1 2
Rser 1 3 0.115
Lser 2 4 0.0000000078
C1 3 4 0.000000012
Rpar 3 4 30000000000
.ends 890334023007_12nF
*******
.subckt 890334023007CS_12nF 1 2
Rser 1 3 0.115
Lser 2 4 0.0000000078
C1 3 4 0.000000012
Rpar 3 4 30000000000
.ends 890334023007CS_12nF
*******
.subckt 890334023008_15nF 1 2
Rser 1 3 0.106
Lser 2 4 0.0000000046
C1 3 4 0.000000015
Rpar 3 4 30000000000
.ends 890334023008_15nF
*******
.subckt 890334023008CS_15nF 1 2
Rser 1 3 0.106
Lser 2 4 0.0000000046
C1 3 4 0.000000015
Rpar 3 4 30000000000
.ends 890334023008CS_15nF
*******
.subckt 890334023010_18nF 1 2
Rser 1 3 0.102
Lser 2 4 0.0000000074
C1 3 4 0.000000018
Rpar 3 4 30000000000
.ends 890334023010_18nF
*******
.subckt 890334023010CS_18nF 1 2
Rser 1 3 0.102
Lser 2 4 0.0000000074
C1 3 4 0.000000018
Rpar 3 4 30000000000
.ends 890334023010CS_18nF
*******
.subckt 890334023011_22nF 1 2
Rser 1 3 0.072
Lser 2 4 0.0000000056
C1 3 4 0.000000022
Rpar 3 4 30000000000
.ends 890334023011_22nF
*******
.subckt 890334023011CS_22nF 1 2
Rser 1 3 0.072
Lser 2 4 0.0000000056
C1 3 4 0.000000022
Rpar 3 4 30000000000
.ends 890334023011CS_22nF
*******
.subckt 890334023015_47nF 1 2
Rser 1 3 0.056
Lser 2 4 0.0000000052
C1 3 4 0.000000047
Rpar 3 4 30000000000
.ends 890334023015_47nF
*******
.subckt 890334023015CS_47nF 1 2
Rser 1 3 0.056
Lser 2 4 0.0000000052
C1 3 4 0.000000047
Rpar 3 4 30000000000
.ends 890334023015CS_47nF
*******
.subckt 890334023017_56nF 1 2
Rser 1 3 0.062
Lser 2 4 0.0000000051
C1 3 4 0.000000056
Rpar 3 4 30000000000
.ends 890334023017_56nF
*******
.subckt 890334023017CS_56nF 1 2
Rser 1 3 0.062
Lser 2 4 0.0000000051
C1 3 4 0.000000056
Rpar 3 4 30000000000
.ends 890334023017CS_56nF
*******
.subckt 890334023019_68nF 1 2
Rser 1 3 0.04
Lser 2 4 0.0000000062
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890334023019_68nF
*******
.subckt 890334023019CS_68nF 1 2
Rser 1 3 0.04
Lser 2 4 0.0000000062
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890334023019CS_68nF
*******
.subckt 890334023021_82nF 1 2
Rser 1 3 0.049
Lser 2 4 0.0000000063
C1 3 4 0.000000082
Rpar 3 4 30000000000
.ends 890334023021_82nF
*******
.subckt 890334023021CS_82nF 1 2
Rser 1 3 0.049
Lser 2 4 0.0000000063
C1 3 4 0.000000082
Rpar 3 4 30000000000
.ends 890334023021CS_82nF
*******
.subckt 890334023023_100nF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000065
C1 3 4 0.0000001
Rpar 3 4 30000000000
.ends 890334023023_100nF
*******
.subckt 890334023023CS_100nF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000065
C1 3 4 0.0000001
Rpar 3 4 30000000000
.ends 890334023023CS_100nF
*******
.subckt 890334023024_120nF 1 2
Rser 1 3 0.043
Lser 2 4 0.0000000057
C1 3 4 0.00000012
Rpar 3 4 30000000000
.ends 890334023024_120nF
*******
.subckt 890334023024CS_120nF 1 2
Rser 1 3 0.043
Lser 2 4 0.0000000057
C1 3 4 0.00000012
Rpar 3 4 30000000000
.ends 890334023024CS_120nF
*******
.subckt 890334023025_150nF 1 2
Rser 1 3 0.045
Lser 2 4 0.0000000056
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890334023025_150nF
*******
.subckt 890334023025CS_150nF 1 2
Rser 1 3 0.045
Lser 2 4 0.0000000056
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890334023025CS_150nF
*******
.subckt 890334023028_220nF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000063
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334023028_220nF
*******
.subckt 890334023028CS_220nF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000063
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334023028CS_220nF
*******
.subckt 890334024001_150nF 1 2
Rser 1 3 0.053
Lser 2 4 0.000000007
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890334024001_150nF
*******
.subckt 890334024001CS_150nF 1 2
Rser 1 3 0.053
Lser 2 4 0.000000007
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890334024001CS_150nF
*******
.subckt 890334024002_220nF 1 2
Rser 1 3 0.043
Lser 2 4 0.00000000586
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334024002_220nF
*******
.subckt 890334024002CS_220nF 1 2
Rser 1 3 0.043
Lser 2 4 0.00000000586
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334024002CS_220nF
*******
.subckt 890334024003_330nF 1 2
Rser 1 3 0.039
Lser 2 4 0.0000000069
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890334024003_330nF
*******
.subckt 890334024003CS_330nF 1 2
Rser 1 3 0.039
Lser 2 4 0.0000000069
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890334024003CS_330nF
*******
.subckt 890334024005_470nF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000068
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890334024005_470nF
*******
.subckt 890334024005CS_470nF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000068
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890334024005CS_470nF
*******
.subckt 890334025004_27nF 1 2
Rser 1 3 0.113
Lser 2 4 0.0000000083
C1 3 4 0.000000027
Rpar 3 4 30000000000
.ends 890334025004_27nF
*******
.subckt 890334025004CS_27nF 1 2
Rser 1 3 0.113
Lser 2 4 0.0000000083
C1 3 4 0.000000027
Rpar 3 4 30000000000
.ends 890334025004CS_27nF
*******
.subckt 890334025006_33nF 1 2
Rser 1 3 0.116
Lser 2 4 0.0000000071
C1 3 4 0.000000033
Rpar 3 4 30000000000
.ends 890334025006_33nF
*******
.subckt 890334025006CS_33nF 1 2
Rser 1 3 0.116
Lser 2 4 0.0000000071
C1 3 4 0.000000033
Rpar 3 4 30000000000
.ends 890334025006CS_33nF
*******
.subckt 890334025007_39nF 1 2
Rser 1 3 0.097
Lser 2 4 0.0000000069
C1 3 4 0.000000039
Rpar 3 4 30000000000
.ends 890334025007_39nF
*******
.subckt 890334025007CS_39nF 1 2
Rser 1 3 0.097
Lser 2 4 0.0000000069
C1 3 4 0.000000039
Rpar 3 4 30000000000
.ends 890334025007CS_39nF
*******
.subckt 890334025009_47nF 1 2
Rser 1 3 0.113
Lser 2 4 0.0000000087
C1 3 4 0.000000047
Rpar 3 4 30000000000
.ends 890334025009_47nF
*******
.subckt 890334025009CS_47nF 1 2
Rser 1 3 0.113
Lser 2 4 0.0000000087
C1 3 4 0.000000047
Rpar 3 4 30000000000
.ends 890334025009CS_47nF
*******
.subckt 890334025011_56nF 1 2
Rser 1 3 0.085
Lser 2 4 0.0000000082
C1 3 4 0.000000056
Rpar 3 4 30000000000
.ends 890334025011_56nF
*******
.subckt 890334025011CS_56nF 1 2
Rser 1 3 0.085
Lser 2 4 0.0000000082
C1 3 4 0.000000056
Rpar 3 4 30000000000
.ends 890334025011CS_56nF
*******
.subckt 890334025013_68nF 1 2
Rser 1 3 0.072
Lser 2 4 0.0000000083
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890334025013_68nF
*******
.subckt 890334025013CS_68nF 1 2
Rser 1 3 0.072
Lser 2 4 0.0000000083
C1 3 4 0.000000068
Rpar 3 4 30000000000
.ends 890334025013CS_68nF
*******
.subckt 890334025015_82nF 1 2
Rser 1 3 0.056
Lser 2 4 0.0000000062
C1 3 4 0.000000082
Rpar 3 4 30000000000
.ends 890334025015_82nF
*******
.subckt 890334025015CS_82nF 1 2
Rser 1 3 0.056
Lser 2 4 0.0000000062
C1 3 4 0.000000082
Rpar 3 4 30000000000
.ends 890334025015CS_82nF
*******
.subckt 890334025017_100nF 1 2
Rser 1 3 0.032
Lser 2 4 0.00000000668
C1 3 4 0.0000001
Rpar 3 4 30000000000
.ends 890334025017_100nF
*******
.subckt 890334025017CS_100nF 1 2
Rser 1 3 0.032
Lser 2 4 0.00000000668
C1 3 4 0.0000001
Rpar 3 4 30000000000
.ends 890334025017CS_100nF
*******
.subckt 890334025020_120nF 1 2
Rser 1 3 0.053
Lser 2 4 0.0000000078
C1 3 4 0.00000012
Rpar 3 4 30000000000
.ends 890334025020_120nF
*******
.subckt 890334025020CS_120nF 1 2
Rser 1 3 0.053
Lser 2 4 0.0000000078
C1 3 4 0.00000012
Rpar 3 4 30000000000
.ends 890334025020CS_120nF
*******
.subckt 890334025022_150nF 1 2
Rser 1 3 0.047
Lser 2 4 0.0000000057
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890334025022_150nF
*******
.subckt 890334025022CS_150nF 1 2
Rser 1 3 0.047
Lser 2 4 0.0000000057
C1 3 4 0.00000015
Rpar 3 4 30000000000
.ends 890334025022CS_150nF
*******
.subckt 890334025025_180nF 1 2
Rser 1 3 0.043
Lser 2 4 0.0000000054
C1 3 4 0.00000018
Rpar 3 4 30000000000
.ends 890334025025_180nF
*******
.subckt 890334025025CS_180nF 1 2
Rser 1 3 0.043
Lser 2 4 0.0000000054
C1 3 4 0.00000018
Rpar 3 4 30000000000
.ends 890334025025CS_180nF
*******
.subckt 890334025027_220nF 1 2
Rser 1 3 0.049
Lser 2 4 0.0000000078
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334025027_220nF
*******
.subckt 890334025027CS_220nF 1 2
Rser 1 3 0.049
Lser 2 4 0.0000000078
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334025027CS_220nF
*******
.subckt 890334025027RP_220nF 1 2
Rser 1 3 0.049
Lser 2 4 0.0000000078
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334025027RP_220nF
*******
.subckt 890334025031_270nF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000091
C1 3 4 0.00000027
Rpar 3 4 30000000000
.ends 890334025031_270nF
*******
.subckt 890334025031CS_270nF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000091
C1 3 4 0.00000027
Rpar 3 4 30000000000
.ends 890334025031CS_270nF
*******
.subckt 890334025034_330nF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000066
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890334025034_330nF
*******
.subckt 890334025034CS_330nF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000066
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890334025034CS_330nF
*******
.subckt 890334025039_470nF 1 2
Rser 1 3 0.037
Lser 2 4 0.0000000065
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890334025039_470nF
*******
.subckt 890334025039CS_470nF 1 2
Rser 1 3 0.037
Lser 2 4 0.0000000065
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890334025039CS_470nF
*******
.subckt 890334025043_560nF 1 2
Rser 1 3 0.027
Lser 2 4 0.0000000072
C1 3 4 0.00000056
Rpar 3 4 17857142857.1429
.ends 890334025043_560nF
*******
.subckt 890334025043CS_560nF 1 2
Rser 1 3 0.027
Lser 2 4 0.0000000072
C1 3 4 0.00000056
Rpar 3 4 17857142857.1429
.ends 890334025043CS_560nF
*******
.subckt 890334025045_680nF 1 2
Rser 1 3 0.027
Lser 2 4 0.0000000085
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890334025045_680nF
*******
.subckt 890334025045CS_680nF 1 2
Rser 1 3 0.027
Lser 2 4 0.0000000085
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890334025045CS_680nF
*******
.subckt 890334026003_220nF 1 2
Rser 1 3 0.061
Lser 2 4 0.00000001323
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334026003_220nF
*******
.subckt 890334026003CS_220nF 1 2
Rser 1 3 0.061
Lser 2 4 0.00000001323
C1 3 4 0.00000022
Rpar 3 4 30000000000
.ends 890334026003CS_220nF
*******
.subckt 890334026007_330nF 1 2
Rser 1 3 0.08
Lser 2 4 0.0000000095
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890334026007_330nF
*******
.subckt 890334026007CS_330nF 1 2
Rser 1 3 0.08
Lser 2 4 0.0000000095
C1 3 4 0.00000033
Rpar 3 4 30000000000
.ends 890334026007CS_330nF
*******
.subckt 890334026014_470nF 1 2
Rser 1 3 0.031
Lser 2 4 0.0000000109
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890334026014_470nF
*******
.subckt 890334026014CS_470nF 1 2
Rser 1 3 0.031
Lser 2 4 0.0000000109
C1 3 4 0.00000047
Rpar 3 4 21276595744.6809
.ends 890334026014CS_470nF
*******
.subckt 890334026018_560nF 1 2
Rser 1 3 0.046
Lser 2 4 0.0000000096
C1 3 4 0.00000056
Rpar 3 4 17857142857.1429
.ends 890334026018_560nF
*******
.subckt 890334026018CS_560nF 1 2
Rser 1 3 0.046
Lser 2 4 0.0000000096
C1 3 4 0.00000056
Rpar 3 4 17857142857.1429
.ends 890334026018CS_560nF
*******
.subckt 890334026020_680nF 1 2
Rser 1 3 0.056
Lser 2 4 0.0000000103
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890334026020_680nF
*******
.subckt 890334026020CS_680nF 1 2
Rser 1 3 0.056
Lser 2 4 0.0000000103
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890334026020CS_680nF
*******
.subckt 890334026024_820nF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000105
C1 3 4 0.00000082
Rpar 3 4 12195121951.2195
.ends 890334026024_820nF
*******
.subckt 890334026024CS_820nF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000105
C1 3 4 0.00000082
Rpar 3 4 12195121951.2195
.ends 890334026024CS_820nF
*******
.subckt 890334026027_1uF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000137
C1 3 4 0.000001
Rpar 3 4 10000000000
.ends 890334026027_1uF
*******
.subckt 890334026027CS_1uF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000137
C1 3 4 0.000001
Rpar 3 4 10000000000
.ends 890334026027CS_1uF
*******
.subckt 890334026030_1.5uF 1 2
Rser 1 3 0.034
Lser 2 4 0.0000000126
C1 3 4 0.0000015
Rpar 3 4 6666666666.66667
.ends 890334026030_1.5uF
*******
.subckt 890334026030CS_1.5uF 1 2
Rser 1 3 0.034
Lser 2 4 0.0000000126
C1 3 4 0.0000015
Rpar 3 4 6666666666.66667
.ends 890334026030CS_1.5uF
*******
.subckt 890334026034_2.2uF 1 2
Rser 1 3 0.025
Lser 2 4 0.0000000105
C1 3 4 0.0000022
Rpar 3 4 4545454545.45455
.ends 890334026034_2.2uF
*******
.subckt 890334026034CS_2.2uF 1 2
Rser 1 3 0.025
Lser 2 4 0.0000000105
C1 3 4 0.0000022
Rpar 3 4 4545454545.45455
.ends 890334026034CS_2.2uF
*******
.subckt 890334027006_680nF 1 2
Rser 1 3 0.035
Lser 2 4 0.0000000135
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890334027006_680nF
*******
.subckt 890334027006CS_680nF 1 2
Rser 1 3 0.035
Lser 2 4 0.0000000135
C1 3 4 0.00000068
Rpar 3 4 14705882352.9412
.ends 890334027006CS_680nF
*******
.subckt 890334027009_1uF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000117
C1 3 4 0.000001
Rpar 3 4 10000000000
.ends 890334027009_1uF
*******
.subckt 890334027009CS_1uF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000117
C1 3 4 0.000001
Rpar 3 4 10000000000
.ends 890334027009CS_1uF
*******
.subckt 890334027012_1.2uF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000168
C1 3 4 0.0000012
Rpar 3 4 8333333333.33333
.ends 890334027012_1.2uF
*******
.subckt 890334027012CS_1.2uF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000168
C1 3 4 0.0000012
Rpar 3 4 8333333333.33333
.ends 890334027012CS_1.2uF
*******
.subckt 890334027021CS_2.2uF 1 2
Rser 1 3 0.019
Lser 2 4 0.000000013
C1 3 4 0.0000022
Rpar 3 4 4545454545.45455
.ends 890334027021CS_2.2uF
*******
.subckt 890334027025_3.3uF 1 2
Rser 1 3 0.023
Lser 2 4 0.0000000139
C1 3 4 0.0000033
Rpar 3 4 3030303030.30303
.ends 890334027025_3.3uF
*******
.subckt 890334027025CS_3.3uF 1 2
Rser 1 3 0.023
Lser 2 4 0.0000000139
C1 3 4 0.0000033
Rpar 3 4 3030303030.30303
.ends 890334027025CS_3.3uF
*******
.subckt 890334027030CS_4.7uF 1 2
Rser 1 3 0.0085
Lser 2 4 0.0000000134
C1 3 4 0.0000047
Rpar 3 4 2127659574.46809
.ends 890334027030CS_4.7uF
*******
.subckt 890334028008_6.8uF 1 2
Rser 1 3 0.015
Lser 2 4 0.0000000135889
C1 3 4 0.0000068
Rpar 3 4 1470588235.29412
.ends 890334028008_6.8uF
*******
.subckt 890334028008CS_6.8uF 1 2
Rser 1 3 0.015
Lser 2 4 0.0000000135889
C1 3 4 0.0000068
Rpar 3 4 1470588235.29412
.ends 890334028008CS_6.8uF
*******
