**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Bi-color Chip LED Waterclear
* Matchcode:              WL-SBCW
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-16
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0606_150066RG74000 1 2 3 4 
D1 4 1 Red
.model Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 3 2 Green
.model Green D
+ IS=75.763E-18
+ N=3.3919
+ RS=.54629
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**************************************************
.subckt 0606_150066SV74000 1 2 3 4
D1 4 1 SRed
.MODEL SRed D
+ IS=17.937E-12
+ N=2.5965
+ RS=.77841
+ IKF=830.60E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 3 2 BGreen
.MODEL BGreen D
+ IS=10.010E-21
+ N=1.9047
+ RS=1.0000E-6
+ IKF=1.0000E3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********************************
.subckt 0606_150066YV74000 1 2 3 4
D1 4 1 Yellow
.MODEL Yellow D
+ IS=6.1031E-15
+ N=2.4355
+ RS=.38909
+ IKF=789.23E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 3 2 BGreen
.MODEL BGreen D
+ IS=15.029E-12
+ N=2.5967
+ RS=.77832
+ IKF=992.81E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********************************
.subckt 1210_150121SV74000 1 2 3 4
D1 4 1 SRed
.MODEL SRed D
+ IS=364.05E-18
+ N=2.2390
+ RS=1.0000E-6
+ IKF=2.1376
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 3 2 BGreen
.MODEL BGreen D
+ IS=10.010E-21
+ N=1.8765
+ RS=1.0000E-6
+ IKF=.18699
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********************************
.subckt 1210_150121YV74000  1 2 3 4
D1 4 1 Yellow
.MODEL Yellow D
+ IS=36.405E-18
+ N=2.2390
+ RS=1.0000E-6
+ IKF=.21375
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 3 2 BGreen
.MODEL BGreen D
+ IS=10.010E-21	
+ N=1.8765
+ RS=1.0000E-6
+ IKF=.18699
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********************************


















