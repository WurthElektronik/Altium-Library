**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  SMT Full-color Chip LED Waterclear
* Matchcode:              WL-SFCW
* Library Type:           LTspice
* Version:                rev22c
* Created/modified by:    Ella      
* Date and Time:          2022-12-14
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0606_150066M173000 1 2 3 4
D1 4 1 Red
.MODEL Red D
+ IS=10.000E-21
+ N=1.7618
+ RS=1.0000E-6
+ IKF=2.0622E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D2 4 2 Green
.MODEL Green D
+ IS=9.0185E-15
+ N=4.0502
+ RS=.65833
+ IKF=796.05E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D3 4 3 Blue 
.MODEL Blue D
+ IS=13.344E-15
+ N=4.1871
+ RS=.69079
+ IKF=802.72E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
.ends
****************************
.subckt 0805_150080M173000 1 2 3 4 
D1 4 1 Red
.MODEL red D
+ IS=10.000E-21
+ N=1.7663
+ RS=1.0000E-6
+ IKF=2.3424E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D2 4 2 Green
.MODEL Green D
+ IS=173.59E-12
+ N=3.9024
+ RS=.92591
+ IKF=155.84E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D3 4 3 Blue 
.MODEL Blue D
+ IS=3.9902E-3
+ N=3.3328
+ RS=.62026
+ IKF=56.277E-18
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
****************************
.subckt 1206_150120M173000 1 2 3 4
D1 2 4 Red
.MODEL Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D2 2 3 Green
.MODEL Green D
+ IS=75.763E-18
+ N=3.3919
+ RS=.54629
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D3 2 1 Blue
.MODEL Blue D
+ IS=48.022E-18
+ N=3.3919
+ RS=.54629
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
****************************
.subckt 1210_150121M173000 1 2 3 4 
D1 4 1 Red
.MODEL Red D
+ IS=10.000E-21
+ N=1.7663
+ RS=1.0004E-6
+ IKF=2.3415E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
D2 4 2 Green
.MODEL Green D
+ IS=3.9902E-3
+ N=3.3328
+ RS=.62026
+ IKF=56.277E-18
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D3 4 3 Blue 
.MODEL Blue D
+ IS=173.59E-12
+ N=3.9024
+ RS=.92591
+ IKF=155.84E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
****************************
.subckt 1206_150120M183000 1 2 3 4
D1 1 2 Red 
.MODEL Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D2 1 3 Blue
.MODEL Blue D
+ IS=48.022E-18
+ N=3.3919
+ RS=.54629
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D3 1 4 Green
.MODEL Green D
+ IS=10.709E-15
+ N=3.2552
+ RS=.77894
+ IKF=7.2378E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
****************************
