**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Infrared Reverse Mount Waterclear Dome
* Matchcode:              WL-SIRW
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-03-01
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1206_15412085A3060 1 2
D1 1 2 SIRW
.MODEL SIRW D
+ IS=10.000E-21
+ N=1.2382
+ RS=1.6930
+ IKF=10.075E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
.ends
*********
.subckt 1206_15412094A3060 1 2
D1 1 2 SIRW
.MODEL SIRW D
+ IS=9.9520E-15
+ N=1.6188
+ RS=.95582
+ IKF=999
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
*********
.subckt 1206_15412085A3060P 1 2
D1 1 2 SIRW
.MODEL SIRW D
+ IS=10.000E-21
+ N=1.2382
+ RS=1.6930
+ IKF=10.075E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*********
.subckt 1206_15412094A3060P 1 2
D1 1 2 SIRW
.MODEL SIRW D
+ IS=9.9520E-15
+ N=1.6188
+ RS=.95582
+ IKF=999
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
*********













































