**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Full-color Chip LED Compact 
* Matchcode:              WL-SFCC
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022/02/16
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0404_150044M155260 1 2 3 4
D1 1 2 Red
.MODEL Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
D2 1 3 Green
.MODEL Green D
+ IS=1.7671E-12
+ N=3.2550
+ RS=.77935
+ IKF=143.59E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
D3 1 4 Blue
.MODEL Blue D
+ IS=829.92E-18
+ N=3.3919
+ RS=.5463
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
.ends
**********
.subckt 0404_150044M155220 1 2 3 4
D1 1 2 Red
.MODEL Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=2.00E-6
+ TT=5.0000E-9
D2 1 3 Blue
.MODEL Blue D
+ IS=270.23E-18
+ N=3.3921
+ RS=.54619
+ IKF=413.52E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=2.00E-6
+ TT=5.0000E-9
D3 1 4 Green
.MODEL Green D
+ IS=237.02E-18
+ N=3.3921
+ RS=.54619
+ IKF=413.52E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=2.00E-6
+ TT=5.0000E-9
.ends
**********