**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT Semi-Shielded Power Inductor
* Matchcode:             WE-LQSA
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         05/31/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
************************************************
.subckt 5040_78404054010_1u 1 2
Rp 1 2 2437
Cp 1 2 1.137p
Rs 1 N3 0.012
L1 N3 2 0.994823u
.ends 5040_78404054010_1u
*******
.subckt 5040_78404054015_1.5u 1 2
Rp 1 2 3015
Cp 1 2 1.325p
Rs 1 N3 0.015
L1 N3 2 1.326u
.ends 5040_78404054015_1.5u
*******
.subckt 5040_78404054022_2.2u 1 2
Rp 1 2 4296
Cp 1 2 3.079p
Rs 1 N3 0.019
L1 N3 2 2.186u
.ends 5040_78404054022_2.2u
*******
.subckt 5040_78404054033_3.3u 1 2
Rp 1 2 5317
Cp 1 2 4.66p
Rs 1 N3 0.024
L1 N3 2 3.233u
.ends 5040_78404054033_3.3u
*******
.subckt 5040_78404054047_4.7u 1 2
Rp 1 2 7273
Cp 1 2 4.297p
Rs 1 N3 0.03
L1 N3 2 4.193u
.ends 5040_78404054047_4.7u
*******
.subckt 5040_78404054068_6.8u 1 2
Rp 1 2 9445
Cp 1 2 4.521p
Rs 1 N3 0.043
L1 N3 2 6.035u
.ends 5040_78404054068_6.8u
*******
.subckt 5040_78404054100_10u 1 2
Rp 1 2 12839
Cp 1 2 4.517p
Rs 1 N3 0.068
L1 N3 2 8.799u
.ends 5040_78404054100_10u
*******
.subckt 5040_78404054150_15u 1 2
Rp 1 2 15690
Cp 1 2 4.916p
Rs 1 N3 0.09
L1 N3 2 13.424u
.ends 5040_78404054150_15u
*******
.subckt 5040_78404054470_47u 1 2
Rp 1 2 28181
Cp 1 2 6.194p
Rs 1 N3 0.29
L1 N3 2 39.832u
.ends 5040_78404054470_47u
*******
.subckt 5040_78404054680_68u 1 2
Rp 1 2 39882
Cp 1 2 5.381p
Rs 1 N3 0.43
L1 N3 2 61.726u
.ends 5040_78404054680_68u
*******
.subckt 5040_78404054101_100u 1 2
Rp 1 2 49818
Cp 1 2 5.441p
Rs 1 N3 0.6
L1 N3 2 89.367u
.ends 5040_78404054101_100u
*******
.subckt 6045_78404064010_1u 1 2
Rp 1 2 2256
Cp 1 2 1.429p
Rs 1 N3 0.009
L1 N3 2 0.791698u
.ends 6045_78404064010_1u
*******
.subckt 6045_78404064015_1.5u 1 2
Rp 1 2 2960
Cp 1 2 1.723p
Rs 1 N3 0.011
L1 N3 2 1.151u
.ends 6045_78404064015_1.5u
*******
.subckt 6045_78404064022_2.2u 1 2
Rp 1 2 4466
Cp 1 2 3.637p
Rs 1 N3 0.014
L1 N3 2 2.071u
.ends 6045_78404064022_2.2u
*******
.subckt 6045_78404064033_3.3u 1 2
Rp 1 2 6090
Cp 1 2 5.476p
Rs 1 N3 0.023
L1 N3 2 3.291u
.ends 6045_78404064033_3.3u
*******
.subckt 6045_78404064047_4.7u 1 2
Rp 1 2 7657
Cp 1 2 5.972p
Rs 1 N3 0.028
L1 N3 2 4.57u
.ends 6045_78404064047_4.7u
*******
.subckt 6045_78404064068_6.8u 1 2
Rp 1 2 8758
Cp 1 2 5.735p
Rs 1 N3 0.035
L1 N3 2 5.822u
.ends 6045_78404064068_6.8u
*******
.subckt 6045_78404064100_10u 1 2
Rp 1 2 11794
Cp 1 2 6.352p
Rs 1 N3 0.048
L1 N3 2 9.034u
.ends 6045_78404064100_10u
*******
.subckt 6045_78404064150_15u 1 2
Rp 1 2 16400
Cp 1 2 7.091p
Rs 1 N3 0.073
L1 N3 2 12.807u
.ends 6045_78404064150_15u
*******
.subckt 6045_78404064220_22u 1 2
Rp 1 2 18664
Cp 1 2 6.566p
Rs 1 N3 0.1
L1 N3 2 18.032u
.ends 6045_78404064220_22u
*******
.subckt 6045_78404064330_33u 1 2
Rp 1 2 26583
Cp 1 2 6.208p
Rs 1 N3 0.14
L1 N3 2 28.912u
.ends 6045_78404064330_33u
*******
.subckt 6045_78404064470_47u 1 2
Rp 1 2 33479
Cp 1 2 6.997p
Rs 1 N3 0.21
L1 N3 2 40.685u
.ends 6045_78404064470_47u
*******
.subckt 6045_78404064680_68u 1 2
Rp 1 2 43031
Cp 1 2 7.379p
Rs 1 N3 0.306
L1 N3 2 61.419u
.ends 6045_78404064680_68u
*******
.subckt 6045_78404064101_100u 1 2
Rp 1 2 43213
Cp 1 2 6.913p
Rs 1 N3 0.443
L1 N3 2 88.257u
.ends 6045_78404064101_100u
*******
.subckt 8040_78404084150_15u 1 2
Rp 1 2 15890
Cp 1 2 5.125p
Rs 1 N3 0.05
L1 N3 2 14.021u
.ends 8040_78404084150_15u
*******
.subckt 8040_78404084220_22u 1 2
Rp 1 2 18454
Cp 1 2 5.956p
Rs 1 N3 0.071
L1 N3 2 19.877u
.ends 8040_78404084220_22u
*******
.subckt 8040_78404084470_33u 1 2
Rp 1 2 30127
Cp 1 2 6.459p
Rs 1 N3 0.14
L1 N3 2 44.077u
.ends 8040_78404084470_33u
*******
.subckt 8040_78404084680_47u 1 2
Rp 1 2 39641
Cp 1 2 6.106p
Rs 1 N3 0.204
L1 N3 2 64.281u
.ends 8040_78404084680_47u
*******
