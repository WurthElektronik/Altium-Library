**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Bi-color Chip LED Compact
* Matchcode:              WL-SBCC
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-09
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0603_150060RV75240 1 2 3 4
D1 3 2 red
.MODEL red D
+ (IS=123.43E-9
+ N=2.5538
+ RS=15.690
+ IKF=14.110E-12
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6)
D2 4 1 bGreen
.MODEL bGreen D
+ (IS=798.77E-12
+ N=4.8320
+ RS=14.210
+ IKF=399.10
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6)
.ends
***********
