**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  MLCCs - Multilayer Ceramic Chip Capacitors
* Matchcode:              WCAP-CSGP_16V
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          07/22/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0201_885012104001_100nF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000008
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0201_885012104001_100nF
*******
.subckt 0201_885012104007_1uF 1 2
Rser 1 3 0.01366
Lser 2 4 0.000000000165
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0201_885012104007_1uF
*******
.subckt 0402_885012005020_1.5pF 1 2
Rser 1 3 1.045
Lser 2 4 0.00000000035
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0402_885012005020_1.5pF
*******
.subckt 0402_885012005021_2.2pF 1 2
Rser 1 3 0.37427104318
Lser 2 4 2.39727122E-10
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0402_885012005021_2.2pF
*******
.subckt 0402_885012005022_3.3pF 1 2
Rser 1 3 0.394048440694
Lser 2 4 2.60787564E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0402_885012005022_3.3pF
*******
.subckt 0402_885012005023_4.7pF 1 2
Rser 1 3 0.475944818481
Lser 2 4 2.97209578E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0402_885012005023_4.7pF
*******
.subckt 0402_885012005024_6.8pF 1 2
Rser 1 3 0.357812051681
Lser 2 4 2.43515953E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0402_885012005024_6.8pF
*******
.subckt 0402_885012005025_10pF 1 2
Rser 1 3 0.486385754904
Lser 2 4 3.42455186E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005025_10pF
*******
.subckt 0402_885012005026_15pF 1 2
Rser 1 3 0.385031326079
Lser 2 4 3.02592165E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885012005026_15pF
*******
.subckt 0402_885012005027_22pF 1 2
Rser 1 3 0.304814718575
Lser 2 4 3.0242914E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885012005027_22pF
*******
.subckt 0402_885012005028_33pF 1 2
Rser 1 3 0.244839252069
Lser 2 4 2.43449082E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005028_33pF
*******
.subckt 0402_885012005029_47pF 1 2
Rser 1 3 0.199232330322
Lser 2 4 2.79396057E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005029_47pF
*******
.subckt 0402_885012005030_68pF 1 2
Rser 1 3 0.183246570883
Lser 2 4 2.43281747E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005030_68pF
*******
.subckt 0402_885012005031_100pF 1 2
Rser 1 3 0.125698815083
Lser 2 4 2.36883012E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005031_100pF
*******
.subckt 0402_885012005032_150pF 1 2
Rser 1 3 0.0914737764723
Lser 2 4 2.04884984E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012005032_150pF
*******
.subckt 0402_885012005033_220pF 1 2
Rser 1 3 0.0784599744138
Lser 2 4 2.05801081E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012005033_220pF
*******
.subckt 0402_885012105014_33nF 1 2
Rser 1 3 0.034439
Lser 2 4 0.000000001077
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0402_885012105014_33nF
*******
.subckt 0402_885012105015_47nF 1 2
Rser 1 3 0.0367849496471
Lser 2 4 1.808767E-10
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0402_885012105015_47nF
*******
.subckt 0402_885012105016_100nF 1 2
Rser 1 3 0.018877276336
Lser 2 4 3.14688963E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012105016_100nF
*******
.subckt 0402_885012105017_220nF 1 2
Rser 1 3 0.0118013539585
Lser 2 4 3.47460059E-10
C1 3 4 0.00000022
Rpar 3 4 500000000
.ends 0402_885012105017_220nF
*******
.subckt 0402_885012205019_100pF 1 2
Rser 1 3 0.77428
Lser 2 4 0.00000000014154
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012205019_100pF
*******
.subckt 0402_885012205020_150pF 1 2
Rser 1 3 0.67192
Lser 2 4 0.00000000015134
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012205020_150pF
*******
.subckt 0402_885012205021_220pF 1 2
Rser 1 3 0.5734
Lser 2 4 0.00000000018579
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012205021_220pF
*******
.subckt 0402_885012205022_330pF 1 2
Rser 1 3 0.41636
Lser 2 4 0.000000000183
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012205022_330pF
*******
.subckt 0402_885012205023_470pF 1 2
Rser 1 3 0.31598
Lser 2 4 0.0000000002154
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012205023_470pF
*******
.subckt 0402_885012205024_680pF 1 2
Rser 1 3 0.23994
Lser 2 4 0.00000000014784
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0402_885012205024_680pF
*******
.subckt 0402_885012205025_1nF 1 2
Rser 1 3 0.213522308242
Lser 2 4 2.15925639E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205025_1nF
*******
.subckt 0402_885012205026_1.5nF 1 2
Rser 1 3 0.17301
Lser 2 4 0.00000000025499
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0402_885012205026_1.5nF
*******
.subckt 0402_885012205027_2.2nF 1 2
Rser 1 3 0.12141
Lser 2 4 0.00000000025109
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0402_885012205027_2.2nF
*******
.subckt 0402_885012205028_3.3nF 1 2
Rser 1 3 0.08715
Lser 2 4 0.00000000022723
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0402_885012205028_3.3nF
*******
.subckt 0402_885012205029_4.7nF 1 2
Rser 1 3 0.07998
Lser 2 4 0.00000000017442
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205029_4.7nF
*******
.subckt 0402_885012205030_6.8nF 1 2
Rser 1 3 0.07283
Lser 2 4 0.00000000019034
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0402_885012205030_6.8nF
*******
.subckt 0402_885012205031_10nF 1 2
Rser 1 3 0.05542
Lser 2 4 0.00000000019893
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0402_885012205031_10nF
*******
.subckt 0402_885012205032_15nF 1 2
Rser 1 3 0.04045
Lser 2 4 0.00000000020744
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0402_885012205032_15nF
*******
.subckt 0402_885012205033_22nF 1 2
Rser 1 3 0.02779
Lser 2 4 0.00000000018757
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0402_885012205033_22nF
*******
.subckt 0402_885012205034_33nF 1 2
Rser 1 3 0.01627
Lser 2 4 0.00000000021013
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0402_885012205034_33nF
*******
.subckt 0402_885012205035_47nF 1 2
Rser 1 3 0.0085
Lser 2 4 0.00000000020707
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0402_885012205035_47nF
*******
.subckt 0402_885012205036_68nF 1 2
Rser 1 3 0.01842
Lser 2 4 0.00000000022333
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0402_885012205036_68nF
*******
.subckt 0402_885012205037_100nF 1 2
Rser 1 3 0.0169137492565
Lser 2 4 3.31963015E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205037_100nF
*******
.subckt 0402_885012205037R_100nF 1 2
Rser 1 3 0.0169137492565
Lser 2 4 3.31963015E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205037R_100nF
*******
.subckt 0402_885012205087_220nF 1 2
Rser 1 3 0.024
Lser 2 4 0.00000000065
C1 3 4 0.00000022
Rpar 3 4 450000000
.ends 0402_885012205087_220nF
*******
.subckt 0402_885012105019_1uF 1 2
Rser 1 3 0.01559
Lser 2 4 0.000000001046
C1 3 4 0.000001
Rpar 3 4 50000000
.ends 0402_885012105019_1uF
*******
.subckt 0603_885012006017_10pF 1 2
Rser 1 3 0.4238423835
Lser 2 4 6.15454653E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006017_10pF
*******
.subckt 0603_885012006018_15pF 1 2
Rser 1 3 0.331903216145
Lser 2 4 4.69540847E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006018_15pF
*******
.subckt 0603_885012006019_22pF 1 2
Rser 1 3 0.348201721723
Lser 2 4 5.50963961E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006019_22pF
*******
.subckt 0603_885012006020_33pF 1 2
Rser 1 3 0.337785757957
Lser 2 4 7.34244223E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006020_33pF
*******
.subckt 0603_885012006021_47pF 1 2
Rser 1 3 0.256261040981
Lser 2 4 6.94150338E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006021_47pF
*******
.subckt 0603_885012006022_68pF 1 2
Rser 1 3 0.161913740901
Lser 2 4 6.38999674E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006022_68pF
*******
.subckt 0603_885012006023_100pF 1 2
Rser 1 3 0.123459009657
Lser 2 4 6.00573816E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006023_100pF
*******
.subckt 0603_885012006024_150pF 1 2
Rser 1 3 0.110788543459
Lser 2 4 5.59777275E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006024_150pF
*******
.subckt 0603_885012006025_220pF 1 2
Rser 1 3 0.0988385216426
Lser 2 4 5.64504761E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012006025_220pF
*******
.subckt 0603_885012006026_330pF 1 2
Rser 1 3 0.0877208643899
Lser 2 4 5.53240043E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006026_330pF
*******
.subckt 0603_885012006027_470pF 1 2
Rser 1 3 0.0602974058901
Lser 2 4 5.48330767E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006027_470pF
*******
.subckt 0603_885012006028_680pF 1 2
Rser 1 3 0.0523826835624
Lser 2 4 5.05789539E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006028_680pF
*******
.subckt 0603_885012006029_1nF 1 2
Rser 1 3 0.0440182000352
Lser 2 4 4.19702079E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006029_1nF
*******
.subckt 0603_885012106013_220nF 1 2
Rser 1 3 0.0111678211386
Lser 2 4 2.40956055E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012106013_220nF
*******
.subckt 0603_885012106014_330nF 1 2
Rser 1 3 0.0117435280097
Lser 2 4 3.10748007E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012106014_330nF
*******
.subckt 0603_885012106015_470nF 1 2
Rser 1 3 0.0117435280097
Lser 2 4 2.50748007E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012106015_470nF
*******
.subckt 0603_885012106016_680nF 1 2
Rser 1 3 0.0127619086118
Lser 2 4 3.65801201E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0603_885012106016_680nF
*******
.subckt 0603_885012106017_1uF 1 2
Rser 1 3 0.00745135412008
Lser 2 4 3.04086627E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012106017_1uF
*******
.subckt 0603_885012106018_2.2uF 1 2
Rser 1 3 0.00721183501635
Lser 2 4 2.59345303E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0603_885012106018_2.2uF
*******
.subckt 0603_885012106029_2.2uF 1 2
Rser 1 3 0.011
Lser 2 4 0.0000000008
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0603_885012106029_2.2uF
*******
.subckt 0603_885012206028_100pF 1 2
Rser 1 3 0.83279
Lser 2 4 0.00000000026283
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206028_100pF
*******
.subckt 0603_885012206029_150pF 1 2
Rser 1 3 0.68443
Lser 2 4 0.00000000029041
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012206029_150pF
*******
.subckt 0603_885012206030_220pF 1 2
Rser 1 3 0.49382
Lser 2 4 0.00000000028774
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012206030_220pF
*******
.subckt 0603_885012206031_330pF 1 2
Rser 1 3 0.4404
Lser 2 4 0.00000000034035
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206031_330pF
*******
.subckt 0603_885012206032_470pF 1 2
Rser 1 3 0.32027
Lser 2 4 0.00000000032279
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206032_470pF
*******
.subckt 0603_885012206033_680pF 1 2
Rser 1 3 0.31076
Lser 2 4 0.00000000037089
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206033_680pF
*******
.subckt 0603_885012206034_1nF 1 2
Rser 1 3 0.2266
Lser 2 4 0.00000000040041
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206034_1nF
*******
.subckt 0603_885012206035_1.5nF 1 2
Rser 1 3 0.13944
Lser 2 4 0.00000000032692
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206035_1.5nF
*******
.subckt 0603_885012206036_2.2nF 1 2
Rser 1 3 0.12185
Lser 2 4 0.00000000030888
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012206036_2.2nF
*******
.subckt 0603_885012206037_3.3nF 1 2
Rser 1 3 0.0993
Lser 2 4 0.00000000030024
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206037_3.3nF
*******
.subckt 0603_885012206038_4.7nF 1 2
Rser 1 3 0.0825557398709
Lser 2 4 2.58966471E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206038_4.7nF
*******
.subckt 0603_885012206039_6.8nF 1 2
Rser 1 3 0.06147
Lser 2 4 0.00000000035083
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206039_6.8nF
*******
.subckt 0603_885012206040_10nF 1 2
Rser 1 3 0.06145
Lser 2 4 0.00000000036058
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206040_10nF
*******
.subckt 0603_885012206041_15nF 1 2
Rser 1 3 0.04438
Lser 2 4 0.00000000031844
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0603_885012206041_15nF
*******
.subckt 0603_885012206042_22nF 1 2
Rser 1 3 0.03181
Lser 2 4 0.00000000024225
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885012206042_22nF
*******
.subckt 0603_885012206043_33nF 1 2
Rser 1 3 0.02195
Lser 2 4 0.00000000030558
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0603_885012206043_33nF
*******
.subckt 0603_885012206044_47nF 1 2
Rser 1 3 0.01525
Lser 2 4 0.00000000027141
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0603_885012206044_47nF
*******
.subckt 0603_885012206045_68nF 1 2
Rser 1 3 0.01508
Lser 2 4 0.00000000030779
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0603_885012206045_68nF
*******
.subckt 0603_885012206046_100nF 1 2
Rser 1 3 0.0189313024822
Lser 2 4 4.50736859E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206046_100nF
*******
.subckt 0603_885012206047_150nF 1 2
Rser 1 3 0.0192205094865
Lser 2 4 4.7670705E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0603_885012206047_150nF
*******
.subckt 0603_885012206048_220nF 1 2
Rser 1 3 0.0139027111992
Lser 2 4 4.40984618E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012206048_220nF
*******
.subckt 0603_885012206049_330nF 1 2
Rser 1 3 0.0117878976558
Lser 2 4 3.9313295E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012206049_330nF
*******
.subckt 0603_885012206050_470nF 1 2
Rser 1 3 0.00930503966198
Lser 2 4 4.27988831E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012206050_470nF
*******
.subckt 0603_885012206051_680nF 1 2
Rser 1 3 0.00730097281816
Lser 2 4 4.2920775E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0603_885012206051_680nF
*******
.subckt 0603_885012206052_1uF 1 2
Rser 1 3 0.00742821402486
Lser 2 4 2.51142993E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0603_885012206052_1uF
*******
.subckt 0805_885012007010_10pF 1 2
Rser 1 3 0.372486331807
Lser 2 4 3.46703717E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0805_885012007010_10pF
*******
.subckt 0805_885012007011_15pF 1 2
Rser 1 3 0.299277635225
Lser 2 4 4.59074821E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007011_15pF
*******
.subckt 0805_885012007012_22pF 1 2
Rser 1 3 0.353164620745
Lser 2 4 4.83956508E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0805_885012007012_22pF
*******
.subckt 0805_885012007013_33pF 1 2
Rser 1 3 0.253567178585
Lser 2 4 4.67181086E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007013_33pF
*******
.subckt 0805_885012007014_47pF 1 2
Rser 1 3 0.224186907869
Lser 2 4 4.55318299E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885012007014_47pF
*******
.subckt 0805_885012007015_68pF 1 2
Rser 1 3 0.177556084991
Lser 2 4 3.40488342E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0805_885012007015_68pF
*******
.subckt 0805_885012007016_100pF 1 2
Rser 1 3 0.144693224126
Lser 2 4 2.25885151E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007016_100pF
*******
.subckt 0805_885012007017_150pF 1 2
Rser 1 3 0.123365902974
Lser 2 4 2.19751744E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007017_150pF
*******
.subckt 0805_885012007018_220pF 1 2
Rser 1 3 0.10837087132
Lser 2 4 2.252525E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012007018_220pF
*******
.subckt 0805_885012007019_330pF 1 2
Rser 1 3 0.0921576071204
Lser 2 4 2.40260993E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007019_330pF
*******
.subckt 0805_885012007020_470pF 1 2
Rser 1 3 0.0750834191209
Lser 2 4 2.93018556E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007020_470pF
*******
.subckt 0805_885012007021_1nF 1 2
Rser 1 3 0.0483999213452
Lser 2 4 2.79211981E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007021_1nF
*******
.subckt 0805_885012007022_1.5nF 1 2
Rser 1 3 0.0373928905809
Lser 2 4 2.95075489E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012007022_1.5nF
*******
.subckt 0805_885012007023_2.2nF 1 2
Rser 1 3 0.0368859488683
Lser 2 4 2.79156194E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012007023_2.2nF
*******
.subckt 0805_885012007024_3.3nF 1 2
Rser 1 3 0.0117602115678
Lser 2 4 2.50664287E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012007024_3.3nF
*******
.subckt 0805_885012007025_4.7nF 1 2
Rser 1 3 0.0198836793746
Lser 2 4 1.51240813E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012007025_4.7nF
*******
.subckt 0805_885012107012_2.2uF 1 2
Rser 1 3 0.0046352610288
Lser 2 4 2.55261723E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012107012_2.2uF
*******
.subckt 0805_885012107013_4.7uF 1 2
Rser 1 3 0.0035599941357
Lser 2 4 2.56410699E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0805_885012107013_4.7uF
*******
.subckt 0805_885012107014_10uF 1 2
Rser 1 3 0.0034022396539
Lser 2 4 3.00259834E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0805_885012107014_10uF
*******
.subckt 0805_885012207027_100pF 1 2
Rser 1 3 0.8158
Lser 2 4 0.00000000024681
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207027_100pF
*******
.subckt 0805_885012207028_150pF 1 2
Rser 1 3 0.69537
Lser 2 4 0.00000000030323
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012207028_150pF
*******
.subckt 0805_885012207029_220pF 1 2
Rser 1 3 0.49653
Lser 2 4 0.00000000027715
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012207029_220pF
*******
.subckt 0805_885012207030_330pF 1 2
Rser 1 3 0.28432
Lser 2 4 0.00000000020282
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012207030_330pF
*******
.subckt 0805_885012207031_470pF 1 2
Rser 1 3 0.19262
Lser 2 4 0.00000000022289
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207031_470pF
*******
.subckt 0805_885012207032_680pF 1 2
Rser 1 3 0.15908
Lser 2 4 0.00000000028074
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012207032_680pF
*******
.subckt 0805_885012207033_1nF 1 2
Rser 1 3 0.10327
Lser 2 4 0.00000000021794
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207033_1nF
*******
.subckt 0805_885012207034_1.5nF 1 2
Rser 1 3 0.0607
Lser 2 4 0.00000000029167
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207034_1.5nF
*******
.subckt 0805_885012207035_2.2nF 1 2
Rser 1 3 0.0294
Lser 2 4 0.00000000027896
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012207035_2.2nF
*******
.subckt 0805_885012207036_3.3nF 1 2
Rser 1 3 0.00336
Lser 2 4 0.00000000024965
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207036_3.3nF
*******
.subckt 0805_885012207037_4.7nF 1 2
Rser 1 3 0.02846
Lser 2 4 0.00000000015236
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012207037_4.7nF
*******
.subckt 0805_885012207038_6.8nF 1 2
Rser 1 3 0.07854
Lser 2 4 0.00000000032137
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0805_885012207038_6.8nF
*******
.subckt 0805_885012207039_10nF 1 2
Rser 1 3 0.06279
Lser 2 4 0.00000000033683
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207039_10nF
*******
.subckt 0805_885012207040_15nF 1 2
Rser 1 3 0.05886
Lser 2 4 0.000000000349367
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0805_885012207040_15nF
*******
.subckt 0805_885012207041_22nF 1 2
Rser 1 3 0.04639
Lser 2 4 0.00000000031523
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0805_885012207041_22nF
*******
.subckt 0805_885012207042_33nF 1 2
Rser 1 3 0.03915
Lser 2 4 0.0000000003028
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0805_885012207042_33nF
*******
.subckt 0805_885012207043_47nF 1 2
Rser 1 3 0.04259
Lser 2 4 0.000000000307
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0805_885012207043_47nF
*******
.subckt 0805_885012207044_68nF 1 2
Rser 1 3 0.02591
Lser 2 4 0.00000000028743
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0805_885012207044_68nF
*******
.subckt 0805_885012207045_100nF 1 2
Rser 1 3 0.0170178433002
Lser 2 4 0.00000000038
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207045_100nF
*******
.subckt 0805_885012207046_150nF 1 2
Rser 1 3 0.0131969599932
Lser 2 4 4.43917137E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0805_885012207046_150nF
*******
.subckt 0805_885012207047_220nF 1 2
Rser 1 3 0.0124886466337
Lser 2 4 0.0000000003
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885012207047_220nF
*******
.subckt 0805_885012207048_330nF 1 2
Rser 1 3 0.0121631731335
Lser 2 4 0.00000000036
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885012207048_330nF
*******
.subckt 0805_885012207049_470nF 1 2
Rser 1 3 0.00820167627427
Lser 2 4 0.00000000049
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0805_885012207049_470nF
*******
.subckt 0805_885012207050_680nF 1 2
Rser 1 3 0.00778029663502
Lser 2 4 0.000000000512
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0805_885012207050_680nF
*******
.subckt 0805_885012207051_1uF 1 2
Rser 1 3 0.0071335712548
Lser 2 4 2.56885128E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885012207051_1uF
*******
.subckt 0805_885012207052_2.2uF 1 2
Rser 1 3 0.00474724521779
Lser 2 4 2.59969084E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012207052_2.2uF
*******
.subckt 0805_885012207053_4.7uF 1 2
Rser 1 3 0.0105
Lser 2 4 0.0000000007
C1 3 4 0.0000047
Rpar 3 4 10000000
.ends 0805_885012207053_4.7uF
*******
.subckt 1206_885012008011_22pF 1 2
Rser 1 3 0.324375840883
Lser 2 4 5.44232375E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1206_885012008011_22pF
*******
.subckt 1206_885012008012_100pF 1 2
Rser 1 3 0.141237836467
Lser 2 4 5.16904289E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008012_100pF
*******
.subckt 1206_885012008013_150pF 1 2
Rser 1 3 0.123922377922
Lser 2 4 4.91328479E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012008013_150pF
*******
.subckt 1206_885012008014_220pF 1 2
Rser 1 3 0.0914487723967
Lser 2 4 4.26746797E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012008014_220pF
*******
.subckt 1206_885012008015_2.2nF 1 2
Rser 1 3 0.0540944991554
Lser 2 4 4.14167967E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012008015_2.2nF
*******
.subckt 1206_885012008016_6.8nF 1 2
Rser 1 3 0.0272311989762
Lser 2 4 3.46260293E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008016_6.8nF
*******
.subckt 1206_885012008017_10nF 1 2
Rser 1 3 0.0157731913832
Lser 2 4 3.49723643E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008017_10nF
*******
.subckt 1206_885012108013_1.5uF 1 2
Rser 1 3 0.0096965404251
Lser 2 4 6.58515557E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 1206_885012108013_1.5uF
*******
.subckt 1206_885012108014_2.2uF 1 2
Rser 1 3 0.00698767716064
Lser 2 4 5.83531315E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012108014_2.2uF
*******
.subckt 1206_885012108015_3.3uF 1 2
Rser 1 3 0.00545085791999
Lser 2 4 6.21772385E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012108015_3.3uF
*******
.subckt 1206_885012108016_4.7uF 1 2
Rser 1 3 0.00700055770575
Lser 2 4 5.37514029E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1206_885012108016_4.7uF
*******
.subckt 1206_885012108017_10uF 1 2
Rser 1 3 0.00377815297038
Lser 2 4 8.77331047E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1206_885012108017_10uF
*******
.subckt 1206_885012108018_22uF 1 2
Rser 1 3 0.00326232270901
Lser 2 4 5.38545474E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1206_885012108018_22uF
*******
.subckt 1206_885012208020_220pF 1 2
Rser 1 3 0.54413
Lser 2 4 0.00000000031019
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012208020_220pF
*******
.subckt 1206_885012208021_470pF 1 2
Rser 1 3 0.34
Lser 2 4 0.00000000042098
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208021_470pF
*******
.subckt 1206_885012208022_1nF 1 2
Rser 1 3 0.23809
Lser 2 4 0.00000000043011
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208022_1nF
*******
.subckt 1206_885012208023_2.2nF 1 2
Rser 1 3 0.16161
Lser 2 4 0.0000000004207
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012208023_2.2nF
*******
.subckt 1206_885012208024_3.3nF 1 2
Rser 1 3 0.12067
Lser 2 4 0.00000000046077
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012208024_3.3nF
*******
.subckt 1206_885012208025_4.7nF 1 2
Rser 1 3 0.1467
Lser 2 4 0.00000000046584
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208025_4.7nF
*******
.subckt 1206_885012208026_10nF 1 2
Rser 1 3 0.07047
Lser 2 4 0.0000000006906
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208026_10nF
*******
.subckt 1206_885012208027_22nF 1 2
Rser 1 3 0.05191
Lser 2 4 0.00000000044884
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1206_885012208027_22nF
*******
.subckt 1206_885012208028_33nF 1 2
Rser 1 3 0.05461
Lser 2 4 0.00000000071542
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1206_885012208028_33nF
*******
.subckt 1206_885012208029_47nF 1 2
Rser 1 3 0.0511
Lser 2 4 0.00000000044681
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1206_885012208029_47nF
*******
.subckt 1206_885012208030_100nF 1 2
Rser 1 3 0.0236394219015
Lser 2 4 6.65660931E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885012208030_100nF
*******
.subckt 1206_885012208031_150nF 1 2
Rser 1 3 0.0172296802581
Lser 2 4 6.75934228E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1206_885012208031_150nF
*******
.subckt 1206_885012208032_220nF 1 2
Rser 1 3 0.0123092011142
Lser 2 4 6.56591189E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1206_885012208032_220nF
*******
.subckt 1206_885012208033_330nF 1 2
Rser 1 3 0.0121092486479
Lser 2 4 7.02655219E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1206_885012208033_330nF
*******
.subckt 1206_885012208034_470nF 1 2
Rser 1 3 0.0106020491014
Lser 2 4 7.42809674E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1206_885012208034_470nF
*******
.subckt 1206_885012208035_680nF 1 2
Rser 1 3 0.00686375950243
Lser 2 4 7.21249479E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1206_885012208035_680nF
*******
.subckt 1206_885012208036_1uF 1 2
Rser 1 3 0.00696547352182
Lser 2 4 6.33927755E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885012208036_1uF
*******
.subckt 1206_885012208037_1.5uF 1 2
Rser 1 3 0.00838199168584
Lser 2 4 6.76254119E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 1206_885012208037_1.5uF
*******
.subckt 1206_885012208038_2.2uF 1 2
Rser 1 3 0.00657322849514
Lser 2 4 5.35127467E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012208038_2.2uF
*******
.subckt 1206_885012208039_3.3uF 1 2
Rser 1 3 0.00583502254442
Lser 2 4 5.58875803E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012208039_3.3uF
*******
.subckt 1206_885012208040_4.7uF 1 2
Rser 1 3 0.00382284206604
Lser 2 4 7.81956777E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1206_885012208040_4.7uF
*******
.subckt 1206_885012208041_10uF 1 2
Rser 1 3 0.00303
Lser 2 4 0.00000000078818
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1206_885012208041_10uF
*******
.subckt 1210_885012009001_15nF 1 2
Rser 1 3 0.0355230024751
Lser 2 4 8.2968558E-11
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1210_885012009001_15nF
*******
.subckt 1210_885012109008_4.7uF 1 2
Rser 1 3 0.0035836083267
Lser 2 4 3.35721238E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012109008_4.7uF
*******
.subckt 1210_885012109009_10uF 1 2
Rser 1 3 0.00244609668461
Lser 2 4 7.73879687E-10
C1 3 4 0.00001
Rpar 3 4 50000000
.ends 1210_885012109009_10uF
*******
.subckt 1210_885012109010_22uF 1 2
Rser 1 3 0.00405759674222
Lser 2 4 1.477484223E-09
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1210_885012109010_22uF
*******
.subckt 1210_885012109011_47uF 1 2
Rser 1 3 0.00321292248127
Lser 2 4 1.005881796E-09
C1 3 4 0.000047
Rpar 3 4 1000000
.ends 1210_885012109011_47uF
*******
.subckt 1210_885012209007_150nF 1 2
Rser 1 3 0.0143454209584
Lser 2 4 5.36188212E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1210_885012209007_150nF
*******
.subckt 1210_885012209008_220nF 1 2
Rser 1 3 0.01034976783
Lser 2 4 5.13522247E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1210_885012209008_220nF
*******
.subckt 1210_885012209009_470nF 1 2
Rser 1 3 0.00837032621271
Lser 2 4 5.45617858E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1210_885012209009_470nF
*******
.subckt 1210_885012209010_680nF 1 2
Rser 1 3 0.00546743874253
Lser 2 4 5.62694253E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1210_885012209010_680nF
*******
.subckt 1210_885012209011_1uF 1 2
Rser 1 3 0.00410122631789
Lser 2 4 3.71398434E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209011_1uF
*******
.subckt 1210_885012209012_2.2uF 1 2
Rser 1 3 0.0039891272832
Lser 2 4 5.25018615E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1210_885012209012_2.2uF
*******
.subckt 1210_885012209013_4.7uF 1 2
Rser 1 3 0.00524566546715
Lser 2 4 5.20085349E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012209013_4.7uF
*******
.subckt 1210_885012209014_10uF 1 2
Rser 1 3 0.00222604043193
Lser 2 4 7.58236705E-10
C1 3 4 0.00001
Rpar 3 4 100000000
.ends 1210_885012209014_10uF
*******
.subckt 1812_885012010001_1nF 1 2
Rser 1 3 0.0510603999373
Lser 2 4 2.97374009E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_885012010001_1nF
*******
.subckt 1812_885012010002_22nF 1 2
Rser 1 3 0.0138901707005
Lser 2 4 3.25297738E-10
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1812_885012010002_22nF
*******
.subckt 1812_885012210001_10nF 1 2
Rser 1 3 0.07465
Lser 2 4 0.00000000052475
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012210001_10nF
*******
.subckt 1812_885012210002_47nF 1 2
Rser 1 3 0.03429
Lser 2 4 0.00000000074448
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1812_885012210002_47nF
*******
.subckt 1812_885012210003_680nF 1 2
Rser 1 3 0.00789799680346
Lser 2 4 5.51300911E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1812_885012210003_680nF
*******
.subckt 1812_885012210004_1uF 1 2
Rser 1 3 0.00726915726357
Lser 2 4 3.95869894E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1812_885012210004_1uF
*******
