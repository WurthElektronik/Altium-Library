**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  SMT Inductor
* Matchcode:              WE-LQ
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Ella
* Date and Time:          12/22/2022
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 1210_744032001_1u  1 2
Rp 1 2 4804.28
Cp 1 2 0.425p
Rs 1 N3 0.08
L1 N3 2 1u
.ends 1210_744032001_1u 
*******
.subckt 1210_7440320015_1.5u  1 2
Rp 1 2 5824.9
Cp 1 2 1.081p
Rs 1 N3 0.104
L1 N3 2 1.5u
.ends 1210_7440320015_1.5u 
*******
.subckt 1210_7440320018_1.8u  1 2
Rp 1 2 6633.9
Cp 1 2 1.494p
Rs 1 N3 0.112
L1 N3 2 1.8u
.ends 1210_7440320018_1.8u 
*******
.subckt 1210_744032002_2.2u  1 2
Rp 1 2 7415.65
Cp 1 2 1.381p
Rs 1 N3 0.12
L1 N3 2 2.2u
.ends 1210_744032002_2.2u 
*******
.subckt 1210_7440320027_2.7u  1 2
Rp 1 2 8345.45
Cp 1 2 1.436p
Rs 1 N3 0.144
L1 N3 2 2.7u
.ends 1210_7440320027_2.7u 
*******
.subckt 1210_744032003_3.3u  1 2
Rp 1 2 10902.3
Cp 1 2 1.338p
Rs 1 N3 0.16
L1 N3 2 3.3u
.ends 1210_744032003_3.3u 
*******
.subckt 1210_7440320039_3.9u  1 2
Rp 1 2 11912.6
Cp 1 2 1.414p
Rs 1 N3 0.2
L1 N3 2 3.9u
.ends 1210_7440320039_3.9u 
*******
.subckt 1210_744032004_4.7u  1 2
Rp 1 2 13116.2
Cp 1 2 1.378p
Rs 1 N3 0.224
L1 N3 2 4.7u
.ends 1210_744032004_4.7u 
*******
.subckt 1210_7440320056_5.6u  1 2
Rp 1 2 15274.5
Cp 1 2 1.258p
Rs 1 N3 0.288
L1 N3 2 5.6u
.ends 1210_7440320056_5.6u 
*******
.subckt 1210_744032006_6.8u  1 2
Rp 1 2 18602.7
Cp 1 2 1.195p
Rs 1 N3 0.32
L1 N3 2 6.8u
.ends 1210_744032006_6.8u 
*******
.subckt 1210_744032008_8.2u  1 2
Rp 1 2 21418.8
Cp 1 2 1.257p
Rs 1 N3 0.36
L1 N3 2 8.2u
.ends 1210_744032008_8.2u 
*******
.subckt 1210_744032100_10u  1 2
Rp 1 2 18455.2
Cp 1 2 1.484p
Rs 1 N3 0.52
L1 N3 2 10u
.ends 1210_744032100_10u 
*******
.subckt 1210_744032101_100u  1 2
Rp 1 2 345196
Cp 1 2 1.985p
Rs 1 N3 5.2
L1 N3 2 100u
.ends 1210_744032101_100u 
*******
.subckt 1210_744032120_12u  1 2
Rp 1 2 26120.9
Cp 1 2 1.56p
Rs 1 N3 0.56
L1 N3 2 12u
.ends 1210_744032120_12u 
*******
.subckt 1210_744032121_120u  1 2
Rp 1 2 91152.9
Cp 1 2 3.805p
Rs 1 N3 5.6
L1 N3 2 120u
.ends 1210_744032121_120u 
*******
.subckt 1210_744032150_15u  1 2
Rp 1 2 30562.4
Cp 1 2 1.391p
Rs 1 N3 0.8
L1 N3 2 15u
.ends 1210_744032150_15u 
*******
.subckt 1210_744032180_18u  1 2
Rp 1 2 32715.2
Cp 1 2 1.555p
Rs 1 N3 0.88
L1 N3 2 18u
.ends 1210_744032180_18u 
*******
.subckt 1210_744032220_22u  1 2
Rp 1 2 30974.7
Cp 1 2 1.677p
Rs 1 N3 1.04
L1 N3 2 22u
.ends 1210_744032220_22u 
*******
.subckt 1210_744032221_220u  1 2
Rp 1 2 1101.39
Cp 1 2 3.355p
Rs 1 N3 9.44
L1 N3 2 220u
.ends 1210_744032221_220u 
*******
.subckt 1210_744032331_330u  1 2
Rp 1 2 389582
Cp 1 2 2.463p
Rs 1 N3 13.2
L1 N3 2 330u
.ends 1210_744032331_330u 
*******
.subckt 1210_744032471_470u  1 2
Rp 1 2 191756
Cp 1 2 5.018p
Rs 1 N3 20
L1 N3 2 470u
.ends 1210_744032471_470u 
*******
.subckt 1210_744032680_68u  1 2
Rp 1 2 63169.1
Cp 1 2 1.883p
Rs 1 N3 3.04
L1 N3 2 68u
.ends 1210_744032680_68u 
*******
.subckt 1210_744032470_47u 1 2
Rp 1 2 63940
Cp 1 2 1.522p
Rs 1 N3 3
L1 N3 2 43.872u
.ends 1210_744032470_47u
*******
.subckt 1812_744045001_1u  1 2
Rp 1 2 4276.73
Cp 1 2 0.424p
Rs 1 N3 0.064
L1 N3 2 1u
.ends 1812_744045001_1u 
*******
.subckt 1812_7440450015_1.5u  1 2
Rp 1 2 3303.93
Cp 1 2 1.155p
Rs 1 N3 0.072
L1 N3 2 1.5u
.ends 1812_7440450015_1.5u 
*******
.subckt 1812_7440450018_1.8u  1 2
Rp 1 2 6268.16
Cp 1 2 0.66p
Rs 1 N3 0.08
L1 N3 2 1.8u
.ends 1812_7440450018_1.8u 
*******
.subckt 1812_744045002_2.2u  1 2
Rp 1 2 7826.16
Cp 1 2 0.863p
Rs 1 N3 0.088
L1 N3 2 2.2u
.ends 1812_744045002_2.2u 
*******
.subckt 1812_7440450027_2.7u  1 2
Rp 1 2 3998.54
Cp 1 2 2.334p
Rs 1 N3 0.096
L1 N3 2 2.7u
.ends 1812_7440450027_2.7u 
*******
.subckt 1812_744045003_3.3u  1 2
Rp 1 2 8748.96
Cp 1 2 2.088p
Rs 1 N3 0.104
L1 N3 2 3.3u
.ends 1812_744045003_3.3u 
*******
.subckt 1812_7440450039_3.9u  1 2
Rp 1 2 10258.6
Cp 1 2 1.976p
Rs 1 N3 0.112
L1 N3 2 3.9u
.ends 1812_7440450039_3.9u 
*******
.subckt 1812_744045004_4.7u  1 2
Rp 1 2 11598.3
Cp 1 2 2.026p
Rs 1 N3 0.12
L1 N3 2 4.7u
.ends 1812_744045004_4.7u 
*******
.subckt 1812_7440450056_5.6u  1 2
Rp 1 2 13756.8
Cp 1 2 1.897p
Rs 1 N3 0.144
L1 N3 2 5.6u
.ends 1812_7440450056_5.6u 
*******
.subckt 1812_744045006_6.8u  1 2
Rp 1 2 13775.2
Cp 1 2 1.988p
Rs 1 N3 0.16
L1 N3 2 6.8u
.ends 1812_744045006_6.8u 
*******
.subckt 1812_744045008_8.2u  1 2
Rp 1 2 15834.6
Cp 1 2 2.012p
Rs 1 N3 0.2
L1 N3 2 8.2u
.ends 1812_744045008_8.2u 
*******
.subckt 1812_744045100_10u  1 2
Rp 1 2 8382.88
Cp 1 2 5.954p
Rs 1 N3 0.24
L1 N3 2 10u
.ends 1812_744045100_10u 
*******
.subckt 1812_744045102_1m  1 2
Rp 1 2 254672
Cp 1 2 4.512p
Rs 1 N3 24
L1 N3 2 1000u
.ends 1812_744045102_1m 
*******
.subckt 1812_744045120_12u  1 2
Rp 1 2 10166.7
Cp 1 2 4.787p
Rs 1 N3 0.336
L1 N3 2 12u
.ends 1812_744045120_12u 
*******
.subckt 1812_744045150_15u  1 2
Rp 1 2 11010.9
Cp 1 2 5.594p
Rs 1 N3 0.4
L1 N3 2 15u
.ends 1812_744045150_15u 
*******
.subckt 1812_744045152_1.5m  1 2
Rp 1 2 280706
Cp 1 2 7.835p
Rs 1 N3 30.8
L1 N3 2 1500u
.ends 1812_744045152_1.5m 
*******
.subckt 1812_744045180_18u  1 2
Rp 1 2 14915.6
Cp 1 2 3.614p
Rs 1 N3 0.48
L1 N3 2 18u
.ends 1812_744045180_18u 
*******
.subckt 1812_744045210_100u  1 2
Rp 1 2 97333.8
Cp 1 2 1.824p
Rs 1 N3 2
L1 N3 2 100u
.ends 1812_744045210_100u 
*******
.subckt 1812_744045215_150u  1 2
Rp 1 2 142715
Cp 1 2 1.852p
Rs 1 N3 2.96
L1 N3 2 150u
.ends 1812_744045215_150u 
*******
.subckt 1812_744045220_22u  1 2
Rp 1 2 33575.6
Cp 1 2 2.229p
Rs 1 N3 0.56
L1 N3 2 22u
.ends 1812_744045220_22u 
*******
.subckt 1812_744045222_2.2m  1 2
Rp 1 2 409779
Cp 1 2 5.677p
Rs 1 N3 50.4
L1 N3 2 2200u
.ends 1812_744045222_2.2m 
*******
.subckt 1812_744045330_33u  1 2
Rp 1 2 44634.5
Cp 1 2 1.74p
Rs 1 N3 0.88
L1 N3 2 33u
.ends 1812_744045330_33u 
*******
.subckt 1812_744045391_390u  1 2
Rp 1 2 125833
Cp 1 2 8.457p
Rs 1 N3 10.4
L1 N3 2 390u
.ends 1812_744045391_390u 
*******
.subckt 1812_744045470_47u  1 2
Rp 1 2 63653
Cp 1 2 2.188p
Rs 1 N3 1.5
L1 N3 2 44.564u
.ends 1812_744045470_47u 
*******
.subckt 1812_744045471_470u  1 2
Rp 1 2 285607
Cp 1 2 3.49p
Rs 1 N3 11.36
L1 N3 2 470u
.ends 1812_744045471_470u 
*******
.subckt 1812_744045681_680u  1 2
Rp 1 2 155713
Cp 1 2 9.454p
Rs 1 N3 13.44
L1 N3 2 680u
.ends 1812_744045681_680u 
*******
.subckt 1812_744045820_82u  1 2
Rp 1 2 176449
Cp 1 2 2.191p
Rs 1 N3 2.3
L1 N3 2 74.804u
.ends 1812_744045820_82u 
*******
.subckt 1812_744045821_820u  1 2
Rp 1 2 165653
Cp 1 2 8.563p
Rs 1 N3 16
L1 N3 2 820u
.ends 1812_744045821_820u 
*******
.subckt 1812_744045680_68u  1 2
Rp 1 2 125000
Cp 1 2 2.2p
Rs 1 N3 2.1
L1 N3 2 60u
.ends 1812_744045680_68u 
*******
