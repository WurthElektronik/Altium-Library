**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Leaded Toroidal Storage Choke
* Matchcode:              WE-SI
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 744101_50u 1 2
Rp 1 2 2496
Cp 1 2 3.228p
Rs 1 N3 0.18
L1 N3 2 50u
.ends 744101_50u
*******
.subckt 744102_73u 1 2
Rp 1 2 3573
Cp 1 2 3.401p
Rs 1 N3 0.23
L1 N3 2 73u
.ends 744102_73u
*******
.subckt 744103_109u 1 2
Rp 1 2 5215
Cp 1 2 4.22p
Rs 1 N3 0.3
L1 N3 2 109u
.ends 744103_109u
*******
.subckt 744104_167u 1 2
Rp 1 2 4827
Cp 1 2 11.727p
Rs 1 N3 0.4
L1 N3 2 167u
.ends 744104_167u
*******
.subckt 744105_258u 1 2
Rp 1 2 6697
Cp 1 2 14.055p
Rs 1 N3 0.4
L1 N3 2 258u
.ends 744105_258u
*******
.subckt 744106_393u 1 2
Rp 1 2 9504
Cp 1 2 16.657p
Rs 1 N3 0.7
L1 N3 2 393u
.ends 744106_393u
*******
.subckt 744107_557u 1 2
Rp 1 2 11007
Cp 1 2 8.991p
Rs 1 N3 0.7
L1 N3 2 557u
.ends 744107_557u
*******
.subckt 744111_37u 1 2
Rp 1 2 1859
Cp 1 2 3.285p
Rs 1 N3 0.6
L1 N3 2 37u
.ends 744111_37u
*******
.subckt 7441110_1.619m 1 2
Rp 1 2 33391
Cp 1 2 52.463p
Rs 1 N3 0.48
L1 N3 2 1886u
.ends 7441110_1.619m
*******
.subckt 744112_53u 1 2
Rp 1 2 2824
Cp 1 2 3.487p
Rs 1 N3 0.8
L1 N3 2 53u
.ends 744112_53u
*******
.subckt 744113_80u 1 2
Rp 1 2 2974
Cp 1 2 10.291p
Rs 1 N3 0.1
L1 N3 2 80u
.ends 744113_80u
*******
.subckt 744114_127u 1 2
Rp 1 2 3286
Cp 1 2 12.89p
Rs 1 N3 0.12
L1 N3 2 127u
.ends 744114_127u
*******
.subckt 744115_200u 1 2
Rp 1 2 5105
Cp 1 2 17.753p
Rs 1 N3 0.2
L1 N3 2 200u
.ends 744115_200u
*******
.subckt 744116_345u 1 2
Rp 1 2 8023
Cp 1 2 27.684p
Rs 1 N3 0.2
L1 N3 2 345u
.ends 744116_345u
*******
.subckt 744117_390u 1 2
Rp 1 2 7419
Cp 1 2 21.675p
Rs 1 N3 0.25
L1 N3 2 390u
.ends 744117_390u
*******
.subckt 744118_600u 1 2
Rp 1 2 11651
Cp 1 2 23.375p
Rs 1 N3 0.33
L1 N3 2 600u
.ends 744118_600u
*******
.subckt 744119_890u 1 2
Rp 1 2 17923
Cp 1 2 37.891p
Rs 1 N3 0.4
L1 N3 2 890u
.ends 744119_890u
*******
.subckt 744131_34u 1 2
Rp 1 2 2079
Cp 1 2 6.846p
Rs 1 N3 0.38
L1 N3 2 34u
.ends 744131_34u
*******
.subckt 744132_49u 1 2
Rp 1 2 2192
Cp 1 2 4.265p
Rs 1 N3 0.5
L1 N3 2 49u
.ends 744132_49u
*******
.subckt 744133_75u 1 2
Rp 1 2 1830
Cp 1 2 4.388p
Rs 1 N3 0.4
L1 N3 2 75u
.ends 744133_75u
*******
.subckt 744134_92u 1 2
Rp 1 2 3470
Cp 1 2 5.871p
Rs 1 N3 0.5
L1 N3 2 92u
.ends 744134_92u
*******
.subckt 744135_157u 1 2
Rp 1 2 4918
Cp 1 2 20.26p
Rs 1 N3 0.63
L1 N3 2 157u
.ends 744135_157u
*******
.subckt 744136_346u 1 2
Rp 1 2 9101
Cp 1 2 8.353p
Rs 1 N3 0.14
L1 N3 2 346u
.ends 744136_346u
*******
.subckt 744137_630u 1 2
Rp 1 2 13135
Cp 1 2 18.884p
Rs 1 N3 0.175
L1 N3 2 630u
.ends 744137_630u
*******
.subckt 744138_727u 1 2
Rp 1 2 12291
Cp 1 2 13.654p
Rs 1 N3 0.24
L1 N3 2 727u
.ends 744138_727u
*******
.subckt 744139_1.124m 1 2
Rp 1 2 22487
Cp 1 2 56.634p
Rs 1 N3 0.28
L1 N3 2 1124u
.ends 744139_1.124m
*******
.subckt 744150_26u 1 2
Rp 1 2 1011
Cp 1 2 4.237p
Rs 1 N3 0.15
L1 N3 2 26u
.ends 744150_26u
*******
.subckt 7441501_12u 1 2
Rp 1 2 629.389
Cp 1 2 1.485p
Rs 1 N3 0.008
L1 N3 2 9.86u
.ends 7441501_12u
*******
.subckt 744151_48u 1 2
Rp 1 2 2470
Cp 1 2 4.961p
Rs 1 N3 0.25
L1 N3 2 48u
.ends 744151_48u
*******
.subckt 744152_82u 1 2
Rp 1 2 2962
Cp 1 2 14.976p
Rs 1 N3 0.3
L1 N3 2 82u
.ends 744152_82u
*******
.subckt 744153_137u 1 2
Rp 1 2 4790
Cp 1 2 7.32p
Rs 1 N3 0.5
L1 N3 2 137u
.ends 744153_137u
*******
.subckt 744154_172u 1 2
Rp 1 2 4572
Cp 1 2 19.529p
Rs 1 N3 0.55
L1 N3 2 172u
.ends 744154_172u
*******
.subckt 744155_220u 1 2
Rp 1 2 3702
Cp 1 2 8.927p
Rs 1 N3 0.6
L1 N3 2 220u
.ends 744155_220u
*******
.subckt 744156_380u 1 2
Rp 1 2 7345
Cp 1 2 33.096p
Rs 1 N3 0.7
L1 N3 2 380u
.ends 744156_380u
*******
