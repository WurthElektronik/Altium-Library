**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Power Inductor 
* Matchcode:              WE-SPC 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 4818_744089410022_0.22u 1 2
Rp 1 2 301.5
Cp 1 2 1.863p
Rs 1 N3 0.015
L1 N3 2 0.22u
.ends 4818_744089410022_0.22u
*******
.subckt 4818_744089410043_0.43u 1 2
Rp 1 2 618.6
Cp 1 2 2.21p
Rs 1 N3 0.0176
L1 N3 2 0.43u
.ends 4818_744089410043_0.43u
*******
.subckt 4818_744089410068_0.68u 1 2
Rp 1 2 980
Cp 1 2 2.635p
Rs 1 N3 0.0221
L1 N3 2 0.68u
.ends 4818_744089410068_0.68u
*******
.subckt 4838_744089430022_0.22u 1 2
Rp 1 2 190
Cp 1 2 0.273p
Rs 1 N3 0.012
L1 N3 2 0.22u
.ends 4838_744089430022_0.22u
*******
.subckt 4838_744089430039_0.39u 1 2
Rp 1 2 310
Cp 1 2 1.8p
Rs 1 N3 0.0135
L1 N3 2 0.39u
.ends 4838_744089430039_0.39u
*******
.subckt 4838_744089430056_0.56u 1 2
Rp 1 2 446
Cp 1 2 2.01p
Rs 1 N3 0.015
L1 N3 2 0.56u
.ends 4838_744089430056_0.56u
*******
.subckt 4838_744089430082_0.82u 1 2
Rp 1 2 700
Cp 1 2 2.28p
Rs 1 N3 0.017
L1 N3 2 0.82u
.ends 4838_744089430082_0.82u
*******
.subckt 4838_74408943010_1u 1 2
Rp 1 2 968
Cp 1 2 2.46p
Rs 1 N3 0.019
L1 N3 2 1u
.ends 4838_74408943010_1u
*******
.subckt 4838_74408943022_2.2u 1 2
Rp 1 2 1820
Cp 1 2 1.65p
Rs 1 N3 0.026
L1 N3 2 2.2u
.ends 4838_74408943022_2.2u
*******
.subckt 4838_74408943033_3.3u 1 2
Rp 1 2 3147
Cp 1 2 3p
Rs 1 N3 0.031
L1 N3 2 3.3u
.ends 4838_74408943033_3.3u
*******
.subckt 4838_74408943047_4.7u 1 2
Rp 1 2 4381
Cp 1 2 3.73p
Rs 1 N3 0.045
L1 N3 2 4.7u
.ends 4838_74408943047_4.7u
*******
.subckt 4838_74408943068_6.8u 1 2
Rp 1 2 6785
Cp 1 2 3.36p
Rs 1 N3 0.051
L1 N3 2 6.8u
.ends 4838_74408943068_6.8u
*******
.subckt 4838_74408943082_8.2u 1 2
Rp 1 2 7275
Cp 1 2 3.7p
Rs 1 N3 0.07
L1 N3 2 8.2u
.ends 4838_74408943082_8.2u
*******
.subckt 4838_74408943100_10u 1 2
Rp 1 2 9380
Cp 1 2 3.24p
Rs 1 N3 0.082
L1 N3 2 10u
.ends 4838_74408943100_10u
*******
.subckt 4838_74408943101_100u 1 2
Rp 1 2 36357
Cp 1 2 6p
Rs 1 N3 0.77
L1 N3 2 100u
.ends 4838_74408943101_100u
*******
.subckt 4838_74408943150_15u 1 2
Rp 1 2 12080
Cp 1 2 3.37p
Rs 1 N3 0.118
L1 N3 2 15u
.ends 4838_74408943150_15u
*******
.subckt 4838_74408943220_22u 1 2
Rp 1 2 17402
Cp 1 2 3.22p
Rs 1 N3 0.185
L1 N3 2 22u
.ends 4838_74408943220_22u
*******
.subckt 4838_74408943330_33u 1 2
Rp 1 2 20970
Cp 1 2 5.54p
Rs 1 N3 0.259
L1 N3 2 33u
.ends 4838_74408943330_33u
*******
.subckt 4838_74408943470_47u 1 2
Rp 1 2 29460
Cp 1 2 5.24p
Rs 1 N3 0.305
L1 N3 2 47u
.ends 4838_74408943470_47u
*******
.subckt 4838_74408943560_56u 1 2
Rp 1 2 22330
Cp 1 2 3.74p
Rs 1 N3 0.418
L1 N3 2 56u
.ends 4838_74408943560_56u
*******
.subckt 4838_74408943680_68u 1 2
Rp 1 2 24666
Cp 1 2 4.48p
Rs 1 N3 0.608
L1 N3 2 68u
.ends 4838_74408943680_68u
*******
.subckt 4838_74408943820_82u 1 2
Rp 1 2 37479
Cp 1 2 5.25p
Rs 1 N3 0.689
L1 N3 2 82u
.ends 4838_74408943820_82u
*******
.subckt 4818_74408941010_1u 1 2
Rp 1 2 1431.9
Cp 1 2 2.79238p
Rs 1 N3 0.0295
L1 N3 2 1u
.ends 4818_74408941010_1u
*******
.subckt 4818_74408941022_2.2u 1 2
Rp 1 2 3588
Cp 1 2 2.76266p
Rs 1 N3 0.06608
L1 N3 2 2.2u
.ends 4818_74408941022_2.2u
*******
.subckt 4818_74408941029_2.9u 1 2
Rp 1 2 4695
Cp 1 2 2.89142p
Rs 1 N3 0.101
L1 N3 2 2.9u
.ends 4818_74408941029_2.9u
*******
.subckt 4818_74408941035_3.5u 1 2
Rp 1 2 5482
Cp 1 2 2.74006p
Rs 1 N3 0.113
L1 N3 2 3.5u
.ends 4818_74408941035_3.5u
*******
.subckt 4818_74408941050_5u 1 2
Rp 1 2 7205
Cp 1 2 2.98886p
Rs 1 N3 0.14
L1 N3 2 5u
.ends 4818_74408941050_5u
*******
.subckt 4818_74408941068_6.8u 1 2
Rp 1 2 10249
Cp 1 2 2.6775p
Rs 1 N3 0.19
L1 N3 2 6.8u
.ends 4818_74408941068_6.8u
*******
.subckt 4818_74408941078_7.8u 1 2
Rp 1 2 11131
Cp 1 2 2.83278p
Rs 1 N3 0.23
L1 N3 2 7.8u
.ends 4818_74408941078_7.8u
*******
.subckt 4818_74408941089_8.9u 1 2
Rp 1 2 12687
Cp 1 2 2.80892p
Rs 1 N3 0.24
L1 N3 2 8.9u
.ends 4818_74408941089_8.9u
*******
.subckt 4818_74408941100_10u 1 2
Rp 1 2 11054
Cp 1 2 2.7239p
Rs 1 N3 0.248
L1 N3 2 10u
.ends 4818_74408941100_10u
*******
.subckt 4818_74408941150_15u 1 2
Rp 1 2 18941
Cp 1 2 3.05924p
Rs 1 N3 0.43
L1 N3 2 15u
.ends 4818_74408941150_15u
*******
.subckt 4818_74408941220_22u 1 2
Rp 1 2 26285
Cp 1 2 3.01946p
Rs 1 N3 0.549
L1 N3 2 22u
.ends 4818_74408941220_22u
*******
.subckt 4818_74408941330_33u 1 2
Rp 1 2 36100
Cp 1 2 3.27186p
Rs 1 N3 1.015
L1 N3 2 33u
.ends 4818_74408941330_33u
*******
.subckt 4818_74408941470_47u 1 2
Rp 1 2 33497
Cp 1 2 2.83752p
Rs 1 N3 1.133
L1 N3 2 47u
.ends 4818_74408941470_47u
*******
.subckt 4828_744089420022_0.22u 1 2
Rp 1 2 244
Cp 1 2 2.11998p
Rs 1 N3 0.0122
L1 N3 2 0.22u
.ends 4828_744089420022_0.22u
*******
.subckt 4828_744089420039_0.39u 1 2
Rp 1 2 427
Cp 1 2 2.35776p
Rs 1 N3 0.015
L1 N3 2 0.39u
.ends 4828_744089420039_0.39u
*******
.subckt 4828_744089420056_0.56u 1 2
Rp 1 2 660
Cp 1 2 2.79788p
Rs 1 N3 0.0156
L1 N3 2 0.56u
.ends 4828_744089420056_0.56u
*******
.subckt 4828_744089420082_0.82u 1 2
Rp 1 2 930
Cp 1 2 2.9594p
Rs 1 N3 0.021
L1 N3 2 0.82u
.ends 4828_744089420082_0.82u
*******
.subckt 4828_74408942012_1.2u 1 2
Rp 1 2 1332
Cp 1 2 3.37718p
Rs 1 N3 0.022
L1 N3 2 1.2u
.ends 4828_74408942012_1.2u
*******
.subckt 4828_74408942022_2.2u 1 2
Rp 1 2 2591
Cp 1 2 3.8222p
Rs 1 N3 0.038
L1 N3 2 2.2u
.ends 4828_74408942022_2.2u
*******
.subckt 4828_74408942033_3.3u 1 2
Rp 1 2 3423
Cp 1 2 4.02904p
Rs 1 N3 0.0483
L1 N3 2 3.3u
.ends 4828_74408942033_3.3u
*******
.subckt 4828_74408942047_4.7u 1 2
Rp 1 2 4627
Cp 1 2 3.70092p
Rs 1 N3 0.0868
L1 N3 2 4.7u
.ends 4828_74408942047_4.7u
*******
.subckt 4828_74408942068_6.8u 1 2
Rp 1 2 5635
Cp 1 2 4.41686p
Rs 1 N3 0.11
L1 N3 2 6.8u
.ends 4828_74408942068_6.8u
*******
.subckt 4828_74408942082_8.2u 1 2
Rp 1 2 6080
Cp 1 2 4.58664p
Rs 1 N3 0.113
L1 N3 2 8.2u
.ends 4828_74408942082_8.2u
*******
.subckt 4828_74408942100_10u 1 2
Rp 1 2 5100
Cp 1 2 4.9144p
Rs 1 N3 0.125
L1 N3 2 10u
.ends 4828_74408942100_10u
*******
.subckt 4828_74408942150_15u 1 2
Rp 1 2 9799
Cp 1 2 4.70946p
Rs 1 N3 0.207
L1 N3 2 15u
.ends 4828_74408942150_15u
*******
.subckt 4828_74408942220_22u 1 2
Rp 1 2 10827
Cp 1 2 5.0532p
Rs 1 N3 0.3
L1 N3 2 22u
.ends 4828_74408942220_22u
*******
.subckt 4828_74408942330_33u 1 2
Rp 1 2 14921
Cp 1 2 5.11808p
Rs 1 N3 0.424
L1 N3 2 33u
.ends 4828_74408942330_33u
*******
.subckt 4828_74408942470_47u 1 2
Rp 1 2 12539
Cp 1 2 6.04294p
Rs 1 N3 0.515
L1 N3 2 47u
.ends 4828_74408942470_47u
*******
.subckt 4828_74408942560_56u 1 2
Rp 1 2 27609
Cp 1 2 5.11108p
Rs 1 N3 0.78
L1 N3 2 56u
.ends 4828_74408942560_56u
*******
.subckt 4828_74408942680_68u 1 2
Rp 1 2 22596
Cp 1 2 6.07534p
Rs 1 N3 0.864
L1 N3 2 68u
.ends 4828_74408942680_68u
*******
.subckt 4828_74408942820_82u 1 2
Rp 1 2 22460
Cp 1 2 5.68162p
Rs 1 N3 0.94
L1 N3 2 82u
.ends 4828_74408942820_82u
*******
