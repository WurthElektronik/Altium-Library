**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Mono-color Ceramic LED Waterclear
* Matchcode:              WL-SMDC
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-21
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 3535_150353BS74500  1  2
D1 1 2  SMDC
.MODEL SMDC D
+ IS=10.000E-21
+ N=2.3829
+ RS=.73019
+ IKF=92.687E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
.ends
******
.subckt 3535_150353GS74500  1  2
D1 1 2 SMDC
.MODEL SMDC D
+ IS=58.235E-18
+ N=3.1569
+ RS=.89951
+ IKF=27.635E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
.ends
******
.subckt 3535_150353RS74500  1  2
D1 1 2 SMDC
.MODEL SMDC D
+ IS=10.000E-21
+ N=1.6253
+ RS=.74692
+ IKF=.10325
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
.ends
******
.subckt 3535_150353YS74500  1  2
D1 1 2 SMDC
.MODEL SMDC D
+ IS=10.000E-21
+ N=1.7107
+ RS=.86724
+ IKF=4.0509
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
.ends
******
.subckt 3535_150353DS74500  1  2
D1 1 2 SMDC
.MODEL SMDC D
+ IS=10.000E-21
+ N=2.3937
+ RS=.70285
+ IKF=98.975E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
.ends
******
.subckt 3535_150353FS74500  1  2
D1 1 2 SMDC
.MODEL SMDC D
+ IS=10.000E-21
+ N=1.4046
+ RS=.45395
+ IKF=79.343E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
.ends
******
.subckt 3535_150353HS74500  1  2
D1 1 2 SMDC
.MODEL SMDC D
+ IS=1.4493E-18
+ N=1.7980
+ RS=1.3215
+ IKF=27.532E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
.ends
******






























































