**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Air Coil 
* Matchcode:              WE-CAIR 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-24
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1322_744910016_1.65n 1 2
C1 1 N7 668.0103f
L1 1 N1 1.5n
L2 N1 N2 23.7775p
L3 N2 N3 61.7144p
L4 N3 N4 313.1481p
L5 N4 N5 78.8413p
L6 N5 N6 56.1893p
R1 2 N1 691.7876m
R2 2 N2 50.7518m
R3 2 N3 31.9165m
R4 2 N4 55.1545m
R5 2 N5 50.9372m
R6 2 N6 59.6202m
R7 2 N7 1.6386
R8 2 1 10g
.ends 
*******
.subckt 1322_744910025_2.55n 1 2
C1 1 N7 724.8882f
L1 1 N1 2.3n
L2 N1 N2 26.4401p
L3 N2 N3 82.2328p
L4 N3 N4 340.1022p
L5 N4 N5 78.9149p
L6 N5 N6 56.2058p
R1 2 N1 685.8509m
R2 2 N2 84.0069m
R3 2 N3 49.3052m
R4 2 N4 55.5305m
R5 2 N5 51.2246m
R6 2 N6 59.8030m
R7 2 N7 1.6452
R8 2 1 10g
.ends 
*******
.subckt 1322_744910038_3.85n 1 2
C1 1 N7 647.8508f
L1 1 N1 3.6n
L2 N1 N2 54.1331p
L3 N2 N3 100.9244p
L4 N3 N4 273.8143p
L5 N4 N5 78.7199p
L6 N5 N6 56.1791p
R1 2 N1 291.6188m
R2 2 N2 93.5354m
R3 2 N3 48.2722m
R4 2 N4 55.0458m
R5 2 N5 51.1528m
R6 2 N6 59.8169m
R7 2 N7 1.631
R8 2 1 10g
.ends 
*******
.subckt 1322_744910054_5.45n 1 2
C1 1 N7 671.4791f
L1 1 N1 5.2n
L2 N1 N2 106.2654p
L3 N2 N3 129.5828p
L4 N3 N4 516.7103p
L5 N4 N5 79.6879p
L6 N5 N6 56.4546p
R1 2 N1 261.4222m
R2 2 N2 134.7785m
R3 2 N3 81.0277m
R4 2 N4 59.9981m
R5 2 N5 55.3527m
R6 2 N6 62.6412m
R7 2 N7 1.6618
R8 2 1 10g
.ends 
*******
.subckt 1340_744911056_5.6n 1 2
C1 1 N7 655.2025f
L1 1 N1 5.4n
L2 N1 N2 127.0466p
L3 N2 N3 135.3291p
L4 N3 N4 154.0151p
L5 N4 N5 177.7449p
L6 N5 N6 156.0717p
R1 2 N1 250.0689m
R2 2 N2 80.8892m
R3 2 N3 56.2504m
R4 2 N4 36.2350m
R5 2 N5 32.7921m
R6 2 N6 48.8656m
R7 2 N7 1.8915
R8 2 1 10g
.ends 
*******
.subckt 1340_744911071_7.15n 1 2
C1 1 N7 655.4814f
L1 1 N1 6.5n
L2 N1 N2 144.1156p
L3 N2 N3 153.5312p
L4 N3 N4 471.7229p
L5 N4 N5 178.8830p
L6 N5 N6 156.2671p
R1 2 N1 262.9679m
R2 2 N2 114.4110m
R3 2 N3 78.4044m
R4 2 N4 46.9462m
R5 2 N5 39.8113m
R6 2 N6 51.2477m
R7 2 N7 1.9952
R8 2 1 10g
.ends 
*******
.subckt 1340_744911088_8.8n 1 2
C1 1 N7 495.4232f
L1 1 N1 8.5n
L2 N1 N2 153.9956p
L3 N2 N3 192.2438p
L4 N3 N4 378.2880p
L5 N4 N5 181.3260p
L6 N5 N6 157.0512p
R1 2 N1 419.1358m
R2 2 N2 168.1055m
R3 2 N3 84.0638m
R4 2 N4 54.4254m
R5 2 N5 49.8872m
R6 2 N6 54.3332m
R7 2 N7 2.5315
R8 2 1 10g
.ends 
*******
.subckt 1340_744911098_9.85n 1 2
C1 1 N7 488.3888f
L1 1 N1 9.5n
L2 N1 N2 202.6653p
L3 N2 N3 247.3084p
L4 N3 N4 1.2288n
L5 N4 N5 185.1519p
L6 N5 N6 158.0064p
R1 2 N1 421.9783m
R2 2 N2 234.4978m
R3 2 N3 155.9979m
R4 2 N4 86.8092m
R5 2 N5 78.5786m
R6 2 N6 76.6357m
R7 2 N7 2.5546
R8 2 1 10g
.ends 
*******
.subckt 1340_744911112_12.55n 1 2
C1 1 N7 347.6595f
L1 1 N1 12n
L2 N1 N2 174.4842p
L3 N2 N3 293.9816p
L4 N3 N4 602.7675p
L5 N4 N5 185.8834p
L6 N5 N6 158.8699p
R1 2 N1 843.4918m
R2 2 N2 270.9034m
R3 2 N3 100.4017m
R4 2 N4 74.9628m
R5 2 N5 71.0115m
R6 2 N6 66.7227m
R7 2 N7 4.4251
R8 2 1 10g
.ends 
*******
.subckt 3136_744913025_2.5n 1 2
C1 1 N7 852.1335f
L1 1 N1 2.3n
L2 N1 N2 38.2717p
L3 N2 N3 637.3483p
L4 N3 N4 755.5919p
L5 N4 N5 178.9546p
L6 N5 N6 156.2103p
R1 2 N1 25.5916m
R2 2 N2 6.2749m
R3 2 N3 25.6713m
R4 2 N4 55.0003m
R5 2 N5 50.6590m
R6 2 N6 59.3872m
R7 2 N7 1.6572
R8 2 1 10g
.ends 
*******
.subckt 3136_744913050_5n 1 2
C1 1 N7 654.0875f
L1 1 N1 4.7n
L2 N1 N2 56.1013p
L3 N2 N3 639.3809p
L4 N3 N4 755.9525p
L5 N4 N5 178.7960p
L6 N5 N6 155.8560p
R1 2 N1 58.9780m
R2 2 N2 19.1272m
R3 2 N3 25.9394m
R4 2 N4 54.9996m
R5 2 N5 50.6518m
R6 2 N6 59.3784m
R7 2 N7 1.6424
R8 2 1 10g
.ends 
*******
.subckt 3136_744913050G_5n 1 2
C1 1 N7 654.0875f
L1 1 N1 4.7n
L2 N1 N2 56.1013p
L3 N2 N3 639.3809p
L4 N3 N4 755.9525p
L5 N4 N5 178.7960p
L6 N5 N6 155.8560p
R1 2 N1 58.9780m
R2 2 N2 19.1272m
R3 2 N3 25.9394m
R4 2 N4 54.9996m
R5 2 N5 50.6518m
R6 2 N6 59.3784m
R7 2 N7 1.6424
R8 2 1 10g
.ends 
*******
.subckt 3136_744913080_8n 1 2
C1 1 N7 550.3851f
L1 1 N1 7.7n
L2 N1 N2 85.4426p
L3 N2 N3 641.4968p
L4 N3 N4 762.6874p
L5 N4 N5 183.8308p
L6 N5 N6 158.9210p
R1 2 N1 117.4271m
R2 2 N2 31.5044m
R3 2 N3 29.7568m
R4 2 N4 55.5761m
R5 2 N5 51.2178m
R6 2 N6 59.7675m
R7 2 N7 2.4173
R8 2 1 10g
.ends 
*******
.subckt 3136_744913080G_8n 1 2
C1 1 N7 550.3851f
L1 1 N1 7.7n
L2 N1 N2 85.4426p
L3 N2 N3 641.4968p
L4 N3 N4 762.6874p
L5 N4 N5 183.8308p
L6 N5 N6 158.9210p
R1 2 N1 117.4271m
R2 2 N2 31.5044m
R3 2 N3 29.7568m
R4 2 N4 55.5761m
R5 2 N5 51.2178m
R6 2 N6 59.7675m
R7 2 N7 2.4173
R8 2 1 10g
.ends 
*******
.subckt 3136_744913112_12.5n 1 2
C1 1 N7 450.9323f
L1 1 N1 12n
L2 N1 N2 116.8776p
L3 N2 N3 682.1951p
L4 N3 N4 795.0749p
L5 N4 N5 199.5531p
L6 N5 N6 163.2640p
R1 2 N1 162.5157m
R2 2 N2 70.6262m
R3 2 N3 97.6940m
R4 2 N4 57.1144m
R5 2 N5 52.4454m
R6 2 N6 60.5189m
R7 2 N7 2.5985
R8 2 1 10g
.ends 
*******
.subckt 3136_744913112G_12.5n 1 2
C1 1 N7 450.9323f
L1 1 N1 12n
L2 N1 N2 116.8776p
L3 N2 N3 682.1951p
L4 N3 N4 795.0749p
L5 N4 N5 199.5531p
L6 N5 N6 163.2640p
R1 2 N1 162.5157m
R2 2 N2 70.6262m
R3 2 N3 97.6940m
R4 2 N4 57.1144m
R5 2 N5 52.4454m
R6 2 N6 60.5189m
R7 2 N7 2.5985
R8 2 1 10g
.ends 
*******
.subckt 3136_744913118_18.5n 1 2
C1 1 N7 512.7156f
L1 1 N1 18n
L2 N1 N2 199.1605p
L3 N2 N3 937.7066p
L4 N3 N4 940.7365p
L5 N4 N5 264.1291p
L6 N5 N6 177.7592p
R1 2 N1 252.6263m
R2 2 N2 108.3958m
R3 2 N3 105.7920m
R4 2 N4 64.7364m
R5 2 N5 58.7177m
R6 2 N6 64.6763m
R7 2 N7 3.292
R8 2 1 10g
.ends 
*******
.subckt 3136_744913118G_18.5n 1 2
C1 1 N7 512.7156f
L1 1 N1 18n
L2 N1 N2 199.1605p
L3 N2 N3 937.7066p
L4 N3 N4 940.7365p
L5 N4 N5 264.1291p
L6 N5 N6 177.7592p
R1 2 N1 252.6263m
R2 2 N2 108.3958m
R3 2 N3 105.7920m
R4 2 N4 64.7364m
R5 2 N5 58.7177m
R6 2 N6 64.6763m
R7 2 N7 3.292
R8 2 1 10g
.ends 
*******
.subckt 3168_744914117_17.5n 1 2
C1 1 N7 202.1713f
L1 1 N1 17n
L2 N1 N2 243.6431p
L3 N2 N3 477.9650p
L4 N3 N4 876.4215p
L5 N4 N5 1.2564n
L6 N5 N6 1.1767n
R1 2 N1 287.2628m
R2 2 N2 72.5845m
R3 2 N3 15.2003m
R4 2 N4 26.5468m
R5 2 N5 38.9202m
R6 2 N6 36.4900m
R7 2 N7 1.436
R8 2 1 10g
.ends 
*******
.subckt 3168_744914117G_17.5n 1 2
C1 1 N7 202.1713f
L1 1 N1 17n
L2 N1 N2 243.6431p
L3 N2 N3 477.9650p
L4 N3 N4 876.4215p
L5 N4 N5 1.2564n
L6 N5 N6 1.1767n
R1 2 N1 287.2628m
R2 2 N2 72.5845m
R3 2 N3 15.2003m
R4 2 N4 26.5468m
R5 2 N5 38.9202m
R6 2 N6 36.4900m
R7 2 N7 1.436
R8 2 1 10g
.ends 
*******
.subckt 3168_744914122_22n 1 2
C1 1 N7 177.0668f
L1 1 N1 21.5n
L2 N1 N2 361.0162p
L3 N2 N3 684.5415p
L4 N3 N4 907.8579p
L5 N4 N5 1.2607n
L6 N5 N6 1.1782n
R1 2 N1 352.9208m
R2 2 N2 80.0586m
R3 2 N3 43.2012m
R4 2 N4 30.9752m
R5 2 N5 39.1554m
R6 2 N6 36.3163m
R7 2 N7 1.6548
R8 2 1 10g
.ends 
*******
.subckt 3168_744914122G_22n 1 2
C1 1 N7 177.0668f
L1 1 N1 21.5n
L2 N1 N2 361.0162p
L3 N2 N3 684.5415p
L4 N3 N4 907.8579p
L5 N4 N5 1.2607n
L6 N5 N6 1.1782n
R1 2 N1 352.9208m
R2 2 N2 80.0586m
R3 2 N3 43.2012m
R4 2 N4 30.9752m
R5 2 N5 39.1554m
R6 2 N6 36.3163m
R7 2 N7 1.6548
R8 2 1 10g
.ends 
*******
.subckt 3168_744914128_28n 1 2
C1 1 N7 176.7787f
L1 1 N1 27.5n
L2 N1 N2 442.0675p
L3 N2 N3 1.2026n
L4 N3 N4 1.0685n
L5 N4 N5 1.3016n
L6 N5 N6 1.1888n
R1 2 N1 464.5980m
R2 2 N2 133.4227m
R3 2 N3 80.7517m
R4 2 N4 53.8611m
R5 2 N5 42.7931m
R6 2 N6 34.9967m
R7 2 N7 2.3901
R8 2 1 10g
.ends 
*******
.subckt 3168_744914128G_28n 1 2
C1 1 N7 176.7787f
L1 1 N1 27.5n
L2 N1 N2 442.0675p
L3 N2 N3 1.2026n
L4 N3 N4 1.0685n
L5 N4 N5 1.3016n
L6 N5 N6 1.1888n
R1 2 N1 464.5980m
R2 2 N2 133.4227m
R3 2 N3 80.7517m
R4 2 N4 53.8611m
R5 2 N5 42.7931m
R6 2 N6 34.9967m
R7 2 N7 2.3901
R8 2 1 10g
.ends 
*******
.subckt 3168_744914135_35.5n 1 2
C1 1 N7 189.0210f
L1 1 N1 35n
L2 N1 N2 603.6856p
L3 N2 N3 1.2544n
L4 N3 N4 1.1156n
L5 N4 N5 1.3267n
L6 N5 N6 1.1956n
R1 2 N1 610.3683m
R2 2 N2 129.6805m
R3 2 N3 84.7788m
R4 2 N4 60.5704m
R5 2 N5 45.8402m
R6 2 N6 34.9666m
R7 2 N7 2.9375
R8 2 1 10g
.ends 
*******
.subckt 3168_744914135G_35.5n 1 2
C1 1 N7 189.0210f
L1 1 N1 35n
L2 N1 N2 603.6856p
L3 N2 N3 1.2544n
L4 N3 N4 1.1156n
L5 N4 N5 1.3267n
L6 N5 N6 1.1956n
R1 2 N1 610.3683m
R2 2 N2 129.6805m
R3 2 N3 84.7788m
R4 2 N4 60.5704m
R5 2 N5 45.8402m
R6 2 N6 34.9666m
R7 2 N7 2.9375
R8 2 1 10g
.ends 
*******
.subckt 3168_744914143_43n 1 2
C1 1 N7 195.1329f
L1 1 N1 42.2n
L2 N1 N2 605.5940p
L3 N2 N3 1.3304n
L4 N3 N4 1.8088n
L5 N4 N5 1.7416n
L6 N5 N6 1.3230n
R1 2 N1 866.7862m
R2 2 N2 214.6286m
R3 2 N3 93.2708m
R4 2 N4 67.7667m
R5 2 N5 49.2671m
R6 2 N6 35.1279m
R7 2 N7 3.1553
R8 2 1 10g
.ends 
*******
.subckt 3168_744914143G_43n 1 2
C1 1 N7 195.1329f
L1 1 N1 42.2n
L2 N1 N2 605.5940p
L3 N2 N3 1.3304n
L4 N3 N4 1.8088n
L5 N4 N5 1.7416n
L6 N5 N6 1.3230n
R1 2 N1 866.7862m
R2 2 N2 214.6286m
R3 2 N3 93.2708m
R4 2 N4 67.7667m
R5 2 N5 49.2671m
R6 2 N6 35.1279m
R7 2 N7 3.1553
R8 2 1 10g
.ends 
*******
.subckt 4248_744912122_22n 1 2
C1 1 N7 176.8930f
L1 1 N1 21.7n
L2 N1 N2 84.3135p
L3 N2 N3 226.3996p
L4 N3 N4 332.2976p
L5 N4 N5 1.6101n
L6 N5 N6 1.3026n
R1 2 N1 479.9697m
R2 2 N2 482.9672m
R3 2 N3 83.7482m
R4 2 N4 66.9750m
R5 2 N5 49.2010m
R6 2 N6 35.2240m
R7 2 N7 3.152
R8 2 1 10g
.ends 
*******
.subckt 4248_744912122G_22n 1 2
C1 1 N7 176.8930f
L1 1 N1 21.7n
L2 N1 N2 84.3135p
L3 N2 N3 226.3996p
L4 N3 N4 332.2976p
L5 N4 N5 1.6101n
L6 N5 N6 1.3026n
R1 2 N1 479.9697m
R2 2 N2 482.9672m
R3 2 N3 83.7482m
R4 2 N4 66.9750m
R5 2 N5 49.2010m
R6 2 N6 35.2240m
R7 2 N7 3.152
R8 2 1 10g
.ends 
*******
.subckt 4248_744912127_27n 1 2
C1 1 N7 215.0029f
L1 1 N1 26.6n
L2 N1 N2 221.1660p
L3 N2 N3 185.5699p
L4 N3 N4 785.2313p
L5 N4 N5 1.5680n
L6 N5 N6 1.3011n
R1 2 N1 471.4079m
R2 2 N2 395.4927m
R3 2 N3 84.9076m
R4 2 N4 66.8938m
R5 2 N5 49.1753m
R6 2 N6 35.2398m
R7 2 N7 2.1629
R8 2 1 10g
.ends 
*******
.subckt 4248_744912127G_27n 1 2
C1 1 N7 215.0029f
L1 1 N1 26.6n
L2 N1 N2 221.1660p
L3 N2 N3 185.5699p
L4 N3 N4 785.2313p
L5 N4 N5 1.5680n
L6 N5 N6 1.3011n
R1 2 N1 471.4079m
R2 2 N2 395.4927m
R3 2 N3 84.9076m
R4 2 N4 66.8938m
R5 2 N5 49.1753m
R6 2 N6 35.2398m
R7 2 N7 2.1629
R8 2 1 10g
.ends 
*******
.subckt 4248_744912133_33n 1 2
C1 1 N7 204.3684f
L1 1 N1 32.5n
L2 N1 N2 263.8048p
L3 N2 N3 268.9599p
L4 N3 N4 830.5381p
L5 N4 N5 1.4260n
L6 N5 N6 1.2920n
R1 2 N1 537.2153m
R2 2 N2 274.5981m
R3 2 N3 87.2485m
R4 2 N4 66.2849m
R5 2 N5 49.0882m
R6 2 N6 35.2747m
R7 2 N7 1.9832
R8 2 1 10g
.ends 
*******
.subckt 4248_744912133G_33n 1 2
C1 1 N7 204.3684f
L1 1 N1 32.5n
L2 N1 N2 263.8048p
L3 N2 N3 268.9599p
L4 N3 N4 830.5381p
L5 N4 N5 1.4260n
L6 N5 N6 1.2920n
R1 2 N1 537.2153m
R2 2 N2 274.5981m
R3 2 N3 87.2485m
R4 2 N4 66.2849m
R5 2 N5 49.0882m
R6 2 N6 35.2747m
R7 2 N7 1.9832
R8 2 1 10g
.ends 
*******
.subckt 4248_744912139_39n 1 2
C1 1 N7 231.9332f
L1 1 N1 38.5n
L2 N1 N2 353.2230p
L3 N2 N3 621.3112p
L4 N3 N4 1.3285n
L5 N4 N5 1.7113n
L6 N5 N6 1.4197n
R1 2 N1 990.9864m
R2 2 N2 210.3492m
R3 2 N3 88.3088m
R4 2 N4 66.6645m
R5 2 N5 49.5817m
R6 2 N6 35.3842m
R7 2 N7 2.1651
R8 2 1 10g
.ends 
*******
.subckt 4248_744912139G_39n 1 2
C1 1 N7 231.9332f
L1 1 N1 38.5n
L2 N1 N2 353.2230p
L3 N2 N3 621.3112p
L4 N3 N4 1.3285n
L5 N4 N5 1.7113n
L6 N5 N6 1.4197n
R1 2 N1 990.9864m
R2 2 N2 210.3492m
R3 2 N3 88.3088m
R4 2 N4 66.6645m
R5 2 N5 49.5817m
R6 2 N6 35.3842m
R7 2 N7 2.1651
R8 2 1 10g
.ends 
*******
.subckt 4248_744912147_47n 1 2
C1 1 N7 244.1549f
L1 1 N1 46.3n
L2 N1 N2 412.9303p
L3 N2 N3 962.9187p
L4 N3 N4 3.9904n
L5 N4 N5 2.5834n
L6 N5 N6 1.6611n
R1 2 N1 1.2043
R2 2 N2 271.6601m
R3 2 N3 101.8974m
R4 2 N4 69.6767m
R5 2 N5 50.3872m
R6 2 N6 34.6274m
R7 2 N7 2.4334
R8 2 1 10g
.ends 
*******
.subckt 4248_744912147G_47n 1 2
C1 1 N7 244.1549f
L1 1 N1 46.3n
L2 N1 N2 412.9303p
L3 N2 N3 962.9187p
L4 N3 N4 3.9904n
L5 N4 N5 2.5834n
L6 N5 N6 1.6611n
R1 2 N1 1.2043
R2 2 N2 271.6601m
R3 2 N3 101.8974m
R4 2 N4 69.6767m
R5 2 N5 50.3872m
R6 2 N6 34.6274m
R7 2 N7 2.4334
R8 2 1 10g
.ends 
*******
.subckt 4248_744912156_56n 1 2
C1 1 N7 272.4250f
L1 1 N1 54n
L2 N1 N2 591.4047p
L3 N2 N3 1.0859n
L4 N3 N4 2.6474n
L5 N4 N5 2.4531n
L6 N5 N6 1.6792n
R1 2 N1 1.4836
R2 2 N2 268.1804m
R3 2 N3 99.5677m
R4 2 N4 67.9343m
R5 2 N5 50.5735m
R6 2 N6 35.1255m
R7 2 N7 2.8276
R8 2 1 10g
.ends 
*******
.subckt 4248_744912156G_56n 1 2
C1 1 N7 272.4250f
L1 1 N1 54n
L2 N1 N2 591.4047p
L3 N2 N3 1.0859n
L4 N3 N4 2.6474n
L5 N4 N5 2.4531n
L6 N5 N6 1.6792n
R1 2 N1 1.4836
R2 2 N2 268.1804m
R3 2 N3 99.5677m
R4 2 N4 67.9343m
R5 2 N5 50.5735m
R6 2 N6 35.1255m
R7 2 N7 2.8276
R8 2 1 10g
.ends 
*******
.subckt 4248_744912168_68n 1 2
C1 1 N7 255.0787f
L1 1 N1 65n
L2 N1 N2 602.0052p
L3 N2 N3 1.1277n
L4 N3 N4 2.6472n
L5 N4 N5 2.4531n
L6 N5 N6 1.6791n
R1 2 N1 1.485
R2 2 N2 274.0530m
R3 2 N3 99.5969m
R4 2 N4 67.9308m
R5 2 N5 50.5730m
R6 2 N6 35.1233m
R7 2 N7 2.828
R8 2 1 10g
.ends 
*******
.subckt 4248_744912168G_68n 1 2
C1 1 N7 255.0787f
L1 1 N1 65n
L2 N1 N2 602.0052p
L3 N2 N3 1.1277n
L4 N3 N4 2.6472n
L5 N4 N5 2.4531n
L6 N5 N6 1.6791n
R1 2 N1 1.485
R2 2 N2 274.0530m
R3 2 N3 99.5969m
R4 2 N4 67.9308m
R5 2 N5 50.5730m
R6 2 N6 35.1233m
R7 2 N7 2.828
R8 2 1 10g
.ends 
*******
.subckt 4248_744912182_82n 1 2
C1 1 N7 305.2065f
L1 1 N1 78n
L2 N1 N2 947.8409p
L3 N2 N3 2.1761n
L4 N3 N4 4.2179n
L5 N4 N5 2.9158n
L6 N5 N6 1.7962n
R1 2 N1 1.5457
R2 2 N2 328.2030m
R3 2 N3 106.2030m
R4 2 N4 70.1066m
R5 2 N5 50.9321m
R6 2 N6 34.4832m
R7 2 N7 2.8371
R8 2 1 10g
.ends 
*******
.subckt 4248_744912182G_82n 1 2
C1 1 N7 305.2065f
L1 1 N1 78n
L2 N1 N2 947.8409p
L3 N2 N3 2.1761n
L4 N3 N4 4.2179n
L5 N4 N5 2.9158n
L6 N5 N6 1.7962n
R1 2 N1 1.5457
R2 2 N2 328.2030m
R3 2 N3 106.2030m
R4 2 N4 70.1066m
R5 2 N5 50.9321m
R6 2 N6 34.4832m
R7 2 N7 2.8371
R8 2 1 10g
.ends 
*******
.subckt 4248_744912210_100n 1 2
C1 1 N7 318.0223f
L1 1 N1 95n
L2 N1 N2 1.1524n
L3 N2 N3 2.4077n
L4 N3 N4 5.7381n
L5 N4 N5 3.4005n
L6 N5 N6 1.9415n
R1 2 N1 1.9587
R2 2 N2 368.6815m
R3 2 N3 118.2784m
R4 2 N4 72.1585m
R5 2 N5 51.1808m
R6 2 N6 33.2519m
R7 2 N7 2.9557
R8 2 1 10g
.ends 
*******
.subckt 4248_744912210G_100n 1 2
C1 1 N7 318.0223f
L1 1 N1 95n
L2 N1 N2 1.1524n
L3 N2 N3 2.4077n
L4 N3 N4 5.7381n
L5 N4 N5 3.4005n
L6 N5 N6 1.9415n
R1 2 N1 1.9587
R2 2 N2 368.6815m
R3 2 N3 118.2784m
R4 2 N4 72.1585m
R5 2 N5 51.1808m
R6 2 N6 33.2519m
R7 2 N7 2.9557
R8 2 1 10g
.ends 
*******
.subckt 4248_744912212_120n 1 2
C1 1 N7 201.7519f
L1 1 N1 115n
L2 N1 N2 1.3134n
L3 N2 N3 2.9094n
L4 N3 N4 6.1371n
L5 N4 N5 3.5035n
L6 N5 N6 1.9755n
R1 2 N1 2.0354
R2 2 N2 405.0626m
R3 2 N3 122.5488m
R4 2 N4 72.7155m
R5 2 N5 51.2271m
R6 2 N6 32.9526m
R7 2 N7 2.9719
R8 2 1 10g
.ends 
*******
.subckt 4248_744912212G_120n 1 2
C1 1 N7 201.7519f
L1 1 N1 115n
L2 N1 N2 1.3134n
L3 N2 N3 2.9094n
L4 N3 N4 6.1371n
L5 N4 N5 3.5035n
L6 N5 N6 1.9755n
R1 2 N1 2.0354
R2 2 N2 405.0626m
R3 2 N3 122.5488m
R4 2 N4 72.7155m
R5 2 N5 51.2271m
R6 2 N6 32.9526m
R7 2 N7 2.9719
R8 2 1 10g
.ends 
*******
.subckt 5910_744918190_90n 1 2
C1 1 N7 385.8930f
L1 1 N1 85.5n
L2 N1 N2 704.1937p
L3 N2 N3 1.4737n
L4 N3 N4 3.4691n
L5 N4 N5 3.0308n
L6 N5 N6 1.9367n
R1 2 N1 1.5246
R2 2 N2 243.0511m
R3 2 N3 77.7824m
R4 2 N4 68.0856m
R5 2 N5 51.6904m
R6 2 N6 35.2838m
R7 2 N7 1.312
R8 2 1 10g
.ends 
*******
.subckt 5910_744918211_111n 1 2
C1 1 N7 352.7334f
L1 1 N1 110n
L2 N1 N2 1.0502n
L3 N2 N3 1.8956n
L4 N3 N4 3.6997n
L5 N4 N5 2.9712n
L6 N5 N6 2.1434n
R1 2 N1 2.59
R2 2 N2 303.2381m
R3 2 N3 112.9595m
R4 2 N4 65.0762m
R5 2 N5 52.3755m
R6 2 N6 35.9450m
R7 2 N7 2.7643
R8 2 1 10g
.ends 
*******
.subckt 5910_744918213_130n 1 2
C1 1 N7 404.6396f
L1 1 N1 128n
L2 N1 N2 1.3366n
L3 N2 N3 2.5222n
L4 N3 N4 5.5807n
L5 N4 N5 3.7075n
L6 N5 N6 2.3592n
R1 2 N1 2.8694
R2 2 N2 348.3838m
R3 2 N3 125.6530m
R4 2 N4 68.3023m
R5 2 N5 53.0464m
R6 2 N6 34.2049m
R7 2 N7 3.3618
R8 2 1 10g
.ends 
*******
.subckt 5910_744918217_169n 1 2
C1 1 N7 372.7053f
L1 1 N1 168n
L2 N1 N2 1.6893n
L3 N2 N3 3.5086n
L4 N3 N4 7.2831n
L5 N4 N5 4.1083n
L6 N5 N6 2.4602n
R1 2 N1 2.9795
R2 2 N2 402.8259m
R3 2 N3 137.9656m
R4 2 N4 71.4227m
R5 2 N5 53.1890m
R6 2 N6 32.7522m
R7 2 N7 3.6178
R8 2 1 10g
.ends 
*******
.subckt 5910_744918220_206n 1 2
C1 1 N7 377.9516f
L1 1 N1 204n
L2 N1 N2 2.1338n
L3 N2 N3 5.2234n
L4 N3 N4 9.1610n
L5 N4 N5 4.4693n
L6 N5 N6 2.5196n
R1 2 N1 3.0851
R2 2 N2 450.6131m
R3 2 N3 152.3304m
R4 2 N4 75.0749m
R5 2 N5 53.0760m
R6 2 N6 30.7841m
R7 2 N7 3.8911
R8 2 1 10g
.ends 
*******
.subckt 5910_744918222_222n 1 2
C1 1 N7 434.6581f
L1 1 N1 218n
L2 N1 N2 2.4014n
L3 N2 N3 5.9031n
L4 N3 N4 10.3234n
L5 N4 N5 4.6760n
L6 N5 N6 2.5380n
R1 2 N1 3.1111
R2 2 N2 517.6863m
R3 2 N3 161.6633m
R4 2 N4 77.3804m
R5 2 N5 52.9011m
R6 2 N6 29.2642m
R7 2 N7 3.9291
R8 2 1 10g
.ends 
*******
.subckt 5910_744918224_246n 1 2
C1 1 N7 420.8593f
L1 1 N1 240n
L2 N1 N2 2.5513n
L3 N2 N3 5.8547n
L4 N3 N4 11.1789n
L5 N4 N5 4.8337n
L6 N5 N6 2.5605n
R1 2 N1 3.1788
R2 2 N2 528.1734m
R3 2 N3 169.7612m
R4 2 N4 79.0638m
R5 2 N5 52.8010m
R6 2 N6 28.0143m
R7 2 N7 4.0104
R8 2 1 10g
.ends 
*******
.subckt 5910_744918230_307n 1 2
C1 1 N7 381.8875f
L1 1 N1 300n
L2 N1 N2 3.3216n
L3 N2 N3 7.7541n
L4 N3 N4 13.8003n
L5 N4 N5 5.1900n
L6 N5 N6 2.5754n
R1 2 N1 3.2722
R2 2 N2 689.3149m
R3 2 N3 202.9174m
R4 2 N4 83.5977m
R5 2 N5 52.5080m
R6 2 N6 24.7691m
R7 2 N7 4.045
R8 2 1 10g
.ends 
*******
.subckt 5910_744918238_380n 1 2
C1 1 N7 394.9573f
L1 1 N1 370n
L2 N1 N2 4.1444n
L3 N2 N3 8.5155n
L4 N3 N4 22.3396n
L5 N4 N5 5.2034n
L6 N5 N6 2.5750n
R1 2 N1 3.2934
R2 2 N2 746.0371m
R3 2 N3 324.6812m
R4 2 N4 83.7697m
R5 2 N5 52.4879m
R6 2 N6 24.5822m
R7 2 N7 4.0588
R8 2 1 10g
.ends 
*******
.subckt 5910_744918242_422n 1 2
C1 1 N7 334.1699f
L1 1 N1 405n
L2 N1 N2 4.8051n
L3 N2 N3 10.5719n
L4 N3 N4 27.3603n
L5 N4 N5 5.2914n
L6 N5 N6 2.6083n
R1 2 N1 3.6452
R2 2 N2 848.6871m
R3 2 N3 396.9749m
R4 2 N4 84.0825m
R5 2 N5 52.6076m
R6 2 N6 24.1782m
R7 2 N7 4.2548
R8 2 1 10g
.ends 
*******
.subckt 5910_744918249_491n 1 2
C1 1 N7 322.6243f
L1 1 N1 470n
L2 N1 N2 5.2373n
L3 N2 N3 17.5130n
L4 N3 N4 40.8475n
L5 N4 N5 6.0813n
L6 N5 N6 3.4447n
R1 2 N1 6.4452
R2 2 N2 868.3077m
R3 2 N3 258.4374m
R4 2 N4 87.5761m
R5 2 N5 56.6037m
R6 2 N6 29.4516m
R7 2 N7 6.5025
R8 2 1 10g
.ends 
*******
.subckt 5910_744918254_538n 1 2
C1 1 N7 365.3684f
L1 1 N1 510n
L2 N1 N2 5.9109n
L3 N2 N3 16.7430n
L4 N3 N4 40.8666n
L5 N4 N5 6.0795n
L6 N5 N6 3.4450n
R1 2 N1 6.4383
R2 2 N2 1.0015
R3 2 N3 284.7418m
R4 2 N4 87.5500m
R5 2 N5 56.6033m
R6 2 N6 29.4596m
R7 2 N7 6.507
R8 2 1 10g
.ends 
*******

