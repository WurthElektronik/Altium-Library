**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ATLL
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 860160272001_22uF 1 2
Rser 1 3 1.70720502503
Lser 2 4 3.491478924E-09
C1 3 4 0.000022
Rpar 3 4 3333333.33333333
.ends 860160272001_22uF
*******
.subckt 860160272002_27uF 1 2
Rser 1 3 1.07993250646
Lser 2 4 3.289117596E-09
C1 3 4 0.000027
Rpar 3 4 3333333.33333333
.ends 860160272002_27uF
*******
.subckt 860160272003_33uF 1 2
Rser 1 3 1.32600426866
Lser 2 4 3.235475421E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860160272003_33uF
*******
.subckt 860160272004_39uF 1 2
Rser 1 3 1.07252972858
Lser 2 4 3.981705347E-09
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860160272004_39uF
*******
.subckt 860160272005_47uF 1 2
Rser 1 3 1.09952414475
Lser 2 4 4.130975975E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860160272005_47uF
*******
.subckt 860160272006_56uF 1 2
Rser 1 3 1.03787598613
Lser 2 4 4.034723783E-09
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860160272006_56uF
*******
.subckt 860160272007_68uF 1 2
Rser 1 3 1.03939605664
Lser 2 4 4.550908878E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860160272007_68uF
*******
.subckt 860160272008_82uF 1 2
Rser 1 3 1.12123323986
Lser 2 4 3.291248461E-09
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860160272008_82uF
*******
.subckt 860160272009_100uF 1 2
Rser 1 3 1.07940871054
Lser 2 4 3.950705111E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860160272009_100uF
*******
.subckt 860160272010_120uF 1 2
Rser 1 3 0.949543169506
Lser 2 4 3.368641777E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860160272010_120uF
*******
.subckt 860160273011_150uF 1 2
Rser 1 3 0.519810933097
Lser 2 4 4.25221849E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860160273011_150uF
*******
.subckt 860160273012_180uF 1 2
Rser 1 3 0.516742077444
Lser 2 4 4.946764876E-09
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160273012_180uF
*******
.subckt 860160273013_220uF 1 2
Rser 1 3 0.33
Lser 2 4 4.231247377E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860160273013_220uF
*******
.subckt 860160273014_270uF 1 2
Rser 1 3 0.305
Lser 2 4 0.0000000028
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860160273014_270uF
*******
.subckt 860160273016_330uF 1 2
Rser 1 3 0.265
Lser 2 4 0.000000003
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160273016_330uF
*******
.subckt 860160273018_390uF 1 2
Rser 1 3 0.195
Lser 2 4 0.000000003
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860160273018_390uF
*******
.subckt 860160273020_470uF 1 2
Rser 1 3 0.233
Lser 2 4 0.0000000029
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860160273020_470uF
*******
.subckt 860160274015_270uF 1 2
Rser 1 3 0.183
Lser 2 4 0.0000000033
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860160274015_270uF
*******
.subckt 860160274017_330uF 1 2
Rser 1 3 0.2
Lser 2 4 0.0000000036
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160274017_330uF
*******
.subckt 860160274019_390uF 1 2
Rser 1 3 0.198
Lser 2 4 0.0000000033
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860160274019_390uF
*******
.subckt 860160274021_470uF 1 2
Rser 1 3 0.206
Lser 2 4 0.0000000032
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860160274021_470uF
*******
.subckt 860160274022_560uF 1 2
Rser 1 3 0.168
Lser 2 4 0.0000000033
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160274022_560uF
*******
.subckt 860160274024_680uF 1 2
Rser 1 3 0.160425711006
Lser 2 4 4.458794028E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860160274024_680uF
*******
.subckt 860160274026_820uF 1 2
Rser 1 3 0.115
Lser 2 4 0.0000000033
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860160274026_820uF
*******
.subckt 860160274029_1mF 1 2
Rser 1 3 0.097
Lser 2 4 0.0000000035
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160274029_1mF
*******
.subckt 860160274032_1.2mF 1 2
Rser 1 3 0.086
Lser 2 4 0.0000000036
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860160274032_1.2mF
*******
.subckt 860160275023_560uF 1 2
Rser 1 3 0.193925509754
Lser 2 4 5.663038306E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160275023_560uF
*******
.subckt 860160275025_680uF 1 2
Rser 1 3 0.121
Lser 2 4 0.0000000042
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860160275025_680uF
*******
.subckt 860160275027_820uF 1 2
Rser 1 3 0.135
Lser 2 4 0.0000000043
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860160275027_820uF
*******
.subckt 860160275028_820uF 1 2
Rser 1 3 0.12622
Lser 2 4 1.2711885515E-08
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860160275028_820uF
*******
.subckt 860160275030_1mF 1 2
Rser 1 3 0.078
Lser 2 4 0.0000000044
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160275030_1mF
*******
.subckt 860160275031_1mF 1 2
Rser 1 3 0.078
Lser 2 4 0.0000000042
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160275031_1mF
*******
.subckt 860160275033_1.2mF 1 2
Rser 1 3 0.082
Lser 2 4 0.0000000037
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860160275033_1.2mF
*******
.subckt 860160275034_1.5mF 1 2
Rser 1 3 0.053
Lser 2 4 0.0000000047
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860160275034_1.5mF
*******
.subckt 860160275035_1.8mF 1 2
Rser 1 3 0.05
Lser 2 4 0.0000000047
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860160275035_1.8mF
*******
.subckt 860160275037_2.2mF 1 2
Rser 1 3 0.041
Lser 2 4 0.0000000042
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860160275037_2.2mF
*******
.subckt 860160275039_2.7mF 1 2
Rser 1 3 0.037
Lser 2 4 0.0000000042
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860160275039_2.7mF
*******
.subckt 860160275041_3.3mF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000044
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860160275041_3.3mF
*******
.subckt 860160278036_1.8mF 1 2
Rser 1 3 0.044
Lser 2 4 0.0000000058
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860160278036_1.8mF
*******
.subckt 860160278038_2.2mF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000054
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860160278038_2.2mF
*******
.subckt 860160278040_2.7mF 1 2
Rser 1 3 0.0441725600168
Lser 2 4 7.882811068E-09
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860160278040_2.7mF
*******
.subckt 860160278042_3.3mF 1 2
Rser 1 3 0.0450086966264
Lser 2 4 8.074795526E-09
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860160278042_3.3mF
*******
.subckt 860160278043_3.9mF 1 2
Rser 1 3 0.0433768094377
Lser 2 4 7.668858814E-09
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860160278043_3.9mF
*******
.subckt 860160278044_4.7mF 1 2
Rser 1 3 0.0363835871313
Lser 2 4 8.311636639E-09
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860160278044_4.7mF
*******
.subckt 860160278046_5.6mF 1 2
Rser 1 3 0.0287918638295
Lser 2 4 7.831495252E-09
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860160278046_5.6mF
*******
.subckt 860160280045_4.7mF 1 2
Rser 1 3 0.0372485963542
Lser 2 4 1.3272088614E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860160280045_4.7mF
*******
.subckt 860160280047_5.6mF 1 2
Rser 1 3 0.0299603444285
Lser 2 4 1.5911637405E-08
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860160280047_5.6mF
*******
.subckt 860160280048_6.8mF 1 2
Rser 1 3 0.0287105349158
Lser 2 4 1.4349391399E-08
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860160280048_6.8mF
*******
.subckt 860160372001_10uF 1 2
Rser 1 3 1.73650604126
Lser 2 4 3.116173958E-09
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 860160372001_10uF
*******
.subckt 860160372002_15uF 1 2
Rser 1 3 1.47774731983
Lser 2 4 3.90470665E-09
C1 3 4 0.000015
Rpar 3 4 5333333.33333333
.ends 860160372002_15uF
*******
.subckt 860160372003_22uF 1 2
Rser 1 3 1.08634572572
Lser 2 4 3.738258747E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860160372003_22uF
*******
.subckt 860160372004_27uF 1 2
Rser 1 3 0.98043238819
Lser 2 4 3.976993288E-09
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 860160372004_27uF
*******
.subckt 860160372005_33uF 1 2
Rser 1 3 1.26947136705
Lser 2 4 5.224380236E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860160372005_33uF
*******
.subckt 860160372006_39uF 1 2
Rser 1 3 1.02212926625
Lser 2 4 3.56775689E-09
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860160372006_39uF
*******
.subckt 860160372007_47uF 1 2
Rser 1 3 0.893291079332
Lser 2 4 4.924322209E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860160372007_47uF
*******
.subckt 860160372008_56uF 1 2
Rser 1 3 0.803469150046
Lser 2 4 4.018347269E-09
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860160372008_56uF
*******
.subckt 860160372009_68uF 1 2
Rser 1 3 0.777295835324
Lser 2 4 4.610268165E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860160372009_68uF
*******
.subckt 860160372011_100uF 1 2
Rser 1 3 0.701709035953
Lser 2 4 3.333375821E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860160372011_100uF
*******
.subckt 860160373010_82uF 1 2
Rser 1 3 0.295
Lser 2 4 0.0000000065
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860160373010_82uF
*******
.subckt 860160373012_120uF 1 2
Rser 1 3 0.3
Lser 2 4 0.0000000029
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860160373012_120uF
*******
.subckt 860160373013_150uF 1 2
Rser 1 3 0.29
Lser 2 4 0.0000000031
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860160373013_150uF
*******
.subckt 860160373014_180uF 1 2
Rser 1 3 0.488703362338
Lser 2 4 4.874044656E-09
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160373014_180uF
*******
.subckt 860160373016_220uF 1 2
Rser 1 3 0.28
Lser 2 4 0.0000000029
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860160373016_220uF
*******
.subckt 860160373018_270uF 1 2
Rser 1 3 0.195
Lser 2 4 0.000000003
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860160373018_270uF
*******
.subckt 860160373021_330uF 1 2
Rser 1 3 0.3088
Lser 2 4 8.200740328E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160373021_330uF
*******
.subckt 860160374015_180uF 1 2
Rser 1 3 0.24
Lser 2 4 0.0000000033
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160374015_180uF
*******
.subckt 860160374017_220uF 1 2
Rser 1 3 0.24
Lser 2 4 0.0000000045
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860160374017_220uF
*******
.subckt 860160374019_270uF 1 2
Rser 1 3 0.21
Lser 2 4 0.0000000032
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860160374019_270uF
*******
.subckt 860160374020_330uF 1 2
Rser 1 3 0.15
Lser 2 4 0.0000000032
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160374020_330uF
*******
.subckt 860160374022_390uF 1 2
Rser 1 3 0.18
Lser 2 4 0.0000000034
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860160374022_390uF
*******
.subckt 860160374024_470uF 1 2
Rser 1 3 0.115
Lser 2 4 0.0000000036
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860160374024_470uF
*******
.subckt 860160374026_560uF 1 2
Rser 1 3 0.09
Lser 2 4 0.0000000035
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160374026_560uF
*******
.subckt 860160374028_680uF 1 2
Rser 1 3 0.139474492952
Lser 2 4 5.279679105E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860160374028_680uF
*******
.subckt 860160374030_820uF 1 2
Rser 1 3 0.063
Lser 2 4 0.0000000035
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860160374030_820uF
*******
.subckt 860160375023_390uF 1 2
Rser 1 3 0.128
Lser 2 4 0.0000000043
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860160375023_390uF
*******
.subckt 860160375025_470uF 1 2
Rser 1 3 0.118
Lser 2 4 0.0000000047
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860160375025_470uF
*******
.subckt 860160375027_560uF 1 2
Rser 1 3 0.152140102566
Lser 2 4 6.241328344E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160375027_560uF
*******
.subckt 860160375029_680uF 1 2
Rser 1 3 0.102564680279
Lser 2 4 4.943659701E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860160375029_680uF
*******
.subckt 860160375031_820uF 1 2
Rser 1 3 0.062
Lser 2 4 0.0000000039
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860160375031_820uF
*******
.subckt 860160375032_1mF 1 2
Rser 1 3 0.058
Lser 2 4 0.000000004
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160375032_1mF
*******
.subckt 860160375033_1.2mF 1 2
Rser 1 3 0.072
Lser 2 4 1.0114544019E-08
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860160375033_1.2mF
*******
.subckt 860160375034_1.5mF 1 2
Rser 1 3 0.045
Lser 2 4 0.0000000046
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860160375034_1.5mF
*******
.subckt 860160375036_1.8mF 1 2
Rser 1 3 0.0487437363971
Lser 2 4 5.509649078E-09
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860160375036_1.8mF
*******
.subckt 860160378035_1.5mF 1 2
Rser 1 3 0.047
Lser 2 4 0.0000000052
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860160378035_1.5mF
*******
.subckt 860160378037_1.8mF 1 2
Rser 1 3 0.041
Lser 2 4 0.0000000056
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860160378037_1.8mF
*******
.subckt 860160378038_2.2mF 1 2
Rser 1 3 0.043
Lser 2 4 0.0000000058
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860160378038_2.2mF
*******
.subckt 860160378039_2.7mF 1 2
Rser 1 3 0.037
Lser 2 4 0.0000000063
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860160378039_2.7mF
*******
.subckt 860160378040_3.3mF 1 2
Rser 1 3 0.0357659071081
Lser 2 4 7.767846599E-09
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860160378040_3.3mF
*******
.subckt 860160378042_3.9mF 1 2
Rser 1 3 0.0308829008546
Lser 2 4 9.49989021E-09
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860160378042_3.9mF
*******
.subckt 860160380041_3.3mF 1 2
Rser 1 3 0.0415014047673
Lser 2 4 1.2758979943E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860160380041_3.3mF
*******
.subckt 860160380043_3.9mF 1 2
Rser 1 3 0.0354654512581
Lser 2 4 1.4845958028E-08
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860160380043_3.9mF
*******
.subckt 860160380044_4.7mF 1 2
Rser 1 3 0.079122135956
Lser 2 4 1.4570249134E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860160380044_4.7mF
*******
.subckt 860160381045_4.7mF 1 2
Rser 1 3 0.0320075532798
Lser 2 4 1.4954913064E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860160381045_4.7mF
*******
.subckt 860160381046_5.6mF 1 2
Rser 1 3 0.0329164494378
Lser 2 4 1.5143018799E-08
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860160381046_5.6mF
*******
.subckt 860160381047_6.8mF 1 2
Rser 1 3 0.0223852751317
Lser 2 4 1.6538948037E-08
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860160381047_6.8mF
*******
.subckt 860160472001_10uF 1 2
Rser 1 3 0.81
Lser 2 4 0.0000000063
C1 3 4 0.00001
Rpar 3 4 8333333.33333333
.ends 860160472001_10uF
*******
.subckt 860160472002_15uF 1 2
Rser 1 3 1.85584013843
Lser 2 4 3.710083353E-09
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends 860160472002_15uF
*******
.subckt 860160472003_22uF 1 2
Rser 1 3 0.773073062777
Lser 2 4 4.185832916E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860160472003_22uF
*******
.subckt 860160472004_27uF 1 2
Rser 1 3 0.964808086736
Lser 2 4 4.67954299E-09
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 860160472004_27uF
*******
.subckt 860160472005_33uF 1 2
Rser 1 3 1.0598402249
Lser 2 4 3.745387003E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860160472005_33uF
*******
.subckt 860160472006_39uF 1 2
Rser 1 3 1.08534229249
Lser 2 4 4.554764183E-09
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860160472006_39uF
*******
.subckt 860160472007_47uF 1 2
Rser 1 3 0.852150045589
Lser 2 4 4.475890707E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860160472007_47uF
*******
.subckt 860160472008_56uF 1 2
Rser 1 3 0.851064971864
Lser 2 4 3.809817688E-09
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860160472008_56uF
*******
.subckt 860160473009_68uF 1 2
Rser 1 3 0.640701805503
Lser 2 4 4.127191313E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860160473009_68uF
*******
.subckt 860160473010_82uF 1 2
Rser 1 3 0.535160810456
Lser 2 4 4.68198713E-09
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860160473010_82uF
*******
.subckt 860160473011_100uF 1 2
Rser 1 3 0.465507875336
Lser 2 4 5.437908885E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860160473011_100uF
*******
.subckt 860160473012_120uF 1 2
Rser 1 3 0.242
Lser 2 4 0.0000000031
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860160473012_120uF
*******
.subckt 860160473013_150uF 1 2
Rser 1 3 0.3
Lser 2 4 0.0000000029
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860160473013_150uF
*******
.subckt 860160473015_180uF 1 2
Rser 1 3 0.248
Lser 2 4 0.000000003
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160473015_180uF
*******
.subckt 860160474014_150uF 1 2
Rser 1 3 0.235
Lser 2 4 0.0000000032
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860160474014_150uF
*******
.subckt 860160474016_180uF 1 2
Rser 1 3 0.17
Lser 2 4 0.0000000034
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160474016_180uF
*******
.subckt 860160474017_220uF 1 2
Rser 1 3 0.15
Lser 2 4 0.0000000033
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860160474017_220uF
*******
.subckt 860160474018_270uF 1 2
Rser 1 3 0.17
Lser 2 4 0.0000000043
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860160474018_270uF
*******
.subckt 860160474019_330uF 1 2
Rser 1 3 0.104
Lser 2 4 0.0000000043
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160474019_330uF
*******
.subckt 860160474021_470uF 1 2
Rser 1 3 0.10968474996
Lser 2 4 4.474658312E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860160474021_470uF
*******
.subckt 860160474023_560uF 1 2
Rser 1 3 0.098
Lser 2 4 0.0000000034
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160474023_560uF
*******
.subckt 860160475020_330uF 1 2
Rser 1 3 0.103
Lser 2 4 0.0000000044
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160475020_330uF
*******
.subckt 860160475022_470uF 1 2
Rser 1 3 0.072
Lser 2 4 0.0000000042
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860160475022_470uF
*******
.subckt 860160475024_560uF 1 2
Rser 1 3 0.077
Lser 2 4 0.0000000042
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160475024_560uF
*******
.subckt 860160475025_680uF 1 2
Rser 1 3 0.061
Lser 2 4 0.0000000046
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860160475025_680uF
*******
.subckt 860160475026_820uF 1 2
Rser 1 3 0.062
Lser 2 4 0.0000000047
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860160475026_820uF
*******
.subckt 860160475027_1mF 1 2
Rser 1 3 0.046
Lser 2 4 0.0000000048
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160475027_1mF
*******
.subckt 860160478028_1mF 1 2
Rser 1 3 0.0665779321447
Lser 2 4 6.593940674E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160478028_1mF
*******
.subckt 860160478029_1.2mF 1 2
Rser 1 3 0.044
Lser 2 4 0.0000000054
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860160478029_1.2mF
*******
.subckt 860160478030_1.5mF 1 2
Rser 1 3 0.0501549106064
Lser 2 4 6.790099498E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860160478030_1.5mF
*******
.subckt 860160478031_1.8mF 1 2
Rser 1 3 0.0372933911506
Lser 2 4 7.773185156E-09
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860160478031_1.8mF
*******
.subckt 860160478033_2.2mF 1 2
Rser 1 3 0.0332489392515
Lser 2 4 8.344397879E-09
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860160478033_2.2mF
*******
.subckt 860160478035_2.7mF 1 2
Rser 1 3 0.0269989842063
Lser 2 4 9.289796954E-09
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860160478035_2.7mF
*******
.subckt 860160480032_1.8mF 1 2
Rser 1 3 0.0397228804443
Lser 2 4 1.3393479845E-08
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860160480032_1.8mF
*******
.subckt 860160480034_2.2mF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000099
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860160480034_2.2mF
*******
.subckt 860160480036_2.7mF 1 2
Rser 1 3 0.0305096809673
Lser 2 4 1.7636663028E-08
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860160480036_2.7mF
*******
.subckt 860160480037_3.3mF 1 2
Rser 1 3 0.0245
Lser 2 4 0.0000000082
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860160480037_3.3mF
*******
.subckt 860160481038_3.3mF 1 2
Rser 1 3 0.0372724932212
Lser 2 4 1.5435087833E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860160481038_3.3mF
*******
.subckt 860160572001_10uF 1 2
Rser 1 3 1.58997939873
Lser 2 4 3.208141074E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860160572001_10uF
*******
.subckt 860160572002_15uF 1 2
Rser 1 3 1.62699209767
Lser 2 4 0.000000003423666
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends 860160572002_15uF
*******
.subckt 860160572003_22uF 1 2
Rser 1 3 1.05275564137
Lser 2 4 3.596801463E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 860160572003_22uF
*******
.subckt 860160572004_27uF 1 2
Rser 1 3 1.15823640158
Lser 2 4 4.2605072E-09
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 860160572004_27uF
*******
.subckt 860160572005_33uF 1 2
Rser 1 3 0.755481675848
Lser 2 4 4.02643178E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860160572005_33uF
*******
.subckt 860160573006_39uF 1 2
Rser 1 3 1.06065726232
Lser 2 4 4.423985835E-09
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860160573006_39uF
*******
.subckt 860160573007_47uF 1 2
Rser 1 3 0.38
Lser 2 4 0.0000000062
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860160573007_47uF
*******
.subckt 860160573008_56uF 1 2
Rser 1 3 0.561017498229
Lser 2 4 5.152586448E-09
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860160573008_56uF
*******
.subckt 860160573009_68uF 1 2
Rser 1 3 0.454317875428
Lser 2 4 3.851305155E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860160573009_68uF
*******
.subckt 860160573010_82uF 1 2
Rser 1 3 0.361240643102
Lser 2 4 5.046495411E-09
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860160573010_82uF
*******
.subckt 860160573012_100uF 1 2
Rser 1 3 327.884758386
Lser 2 4 4.790890144E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860160573012_100uF
*******
.subckt 860160574011_82uF 1 2
Rser 1 3 0.18
Lser 2 4 0.0000000078
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860160574011_82uF
*******
.subckt 860160574013_100uF 1 2
Rser 1 3 0.18
Lser 2 4 0.0000000033
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860160574013_100uF
*******
.subckt 860160574014_120uF 1 2
Rser 1 3 0.16
Lser 2 4 0.0000000033
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860160574014_120uF
*******
.subckt 860160574015_150uF 1 2
Rser 1 3 0.18
Lser 2 4 0.000000003
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860160574015_150uF
*******
.subckt 860160574017_180uF 1 2
Rser 1 3 0.143
Lser 2 4 0.0000000034
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160574017_180uF
*******
.subckt 860160574019_220uF 1 2
Rser 1 3 0.128
Lser 2 4 0.0000000035
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860160574019_220uF
*******
.subckt 860160574021_270uF 1 2
Rser 1 3 0.105
Lser 2 4 0.0000000032
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860160574021_270uF
*******
.subckt 860160574023_330uF 1 2
Rser 1 3 0.083
Lser 2 4 0.0000000032
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160574023_330uF
*******
.subckt 860160575016_150uF 1 2
Rser 1 3 0.224289676301
Lser 2 4 5.241169216E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860160575016_150uF
*******
.subckt 860160575018_180uF 1 2
Rser 1 3 0.155
Lser 2 4 0.0000000046
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160575018_180uF
*******
.subckt 860160575020_220uF 1 2
Rser 1 3 0.156026739829
Lser 2 4 7.35923697E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860160575020_220uF
*******
.subckt 860160575022_270uF 1 2
Rser 1 3 0.169121030463
Lser 2 4 7.290579128E-09
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860160575022_270uF
*******
.subckt 860160575024_330uF 1 2
Rser 1 3 0.0966735056039
Lser 2 4 5.188451025E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160575024_330uF
*******
.subckt 860160575025_470uF 1 2
Rser 1 3 0.067
Lser 2 4 0.0000000049
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860160575025_470uF
*******
.subckt 860160575026_560uF 1 2
Rser 1 3 0.0699097504914
Lser 2 4 5.682141396E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160575026_560uF
*******
.subckt 860160575028_680uF 1 2
Rser 1 3 0.058
Lser 2 4 0.0000000047
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860160575028_680uF
*******
.subckt 860160575031_1mF 1 2
Rser 1 3 0.0377413960237
Lser 2 4 5.417475882E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160575031_1mF
*******
.subckt 860160578027_560uF 1 2
Rser 1 3 0.051
Lser 2 4 0.0000000057
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160578027_560uF
*******
.subckt 860160578029_680uF 1 2
Rser 1 3 0.046
Lser 2 4 0.0000000055
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860160578029_680uF
*******
.subckt 860160578030_820uF 1 2
Rser 1 3 0.0517134439344
Lser 2 4 6.329298467E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860160578030_820uF
*******
.subckt 860160578032_1mF 1 2
Rser 1 3 0.0348198334666
Lser 2 4 8.331084265E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160578032_1mF
*******
.subckt 860160578033_1.2mF 1 2
Rser 1 3 0.040908356763
Lser 2 4 7.297550453E-09
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860160578033_1.2mF
*******
.subckt 860160578034_1.5mF 1 2
Rser 1 3 0.0267010589013
Lser 2 4 9.006874728E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860160578034_1.5mF
*******
.subckt 860160578036_1.8mF 1 2
Rser 1 3 0.0277173048429
Lser 2 4 8.996635861E-09
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860160578036_1.8mF
*******
.subckt 860160580035_1.5mF 1 2
Rser 1 3 0.026
Lser 2 4 0.0000000075
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860160580035_1.5mF
*******
.subckt 860160580037_1.8mF 1 2
Rser 1 3 0.0313464987027
Lser 2 4 1.5813035608E-08
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860160580037_1.8mF
*******
.subckt 860160580038_2.2mF 1 2
Rser 1 3 0.0273252373753
Lser 2 4 1.3391011252E-08
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860160580038_2.2mF
*******
.subckt 860160581039_2.2mF 1 2
Rser 1 3 0.0329576211809
Lser 2 4 1.5018684306E-08
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860160581039_2.2mF
*******
.subckt 860160581040_2.7mF 1 2
Rser 1 3 0.0271774285032
Lser 2 4 1.4703601729E-08
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860160581040_2.7mF
*******
.subckt 860160672001_470nF 1 2
Rser 1 3 2.33587961101
Lser 2 4 2.335951402E-09
C1 3 4 0.00000047
Rpar 3 4 16666666.6666667
.ends 860160672001_470nF
*******
.subckt 860160672002_1uF 1 2
Rser 1 3 2.22482284088
Lser 2 4 3.144700229E-09
C1 3 4 0.000001
Rpar 3 4 16666666.6666667
.ends 860160672002_1uF
*******
.subckt 860160672003_2.2uF 1 2
Rser 1 3 0.92
Lser 2 4 0.000000005
C1 3 4 0.0000022
Rpar 3 4 16666666.6666667
.ends 860160672003_2.2uF
*******
.subckt 860160672004_3.3uF 1 2
Rser 1 3 1.23768720729
Lser 2 4 3.712648854E-09
C1 3 4 0.0000033
Rpar 3 4 16666666.6666667
.ends 860160672004_3.3uF
*******
.subckt 860160672005_4.7uF 1 2
Rser 1 3 1.68223154882
Lser 2 4 3.143769413E-09
C1 3 4 0.0000047
Rpar 3 4 16666666.6666667
.ends 860160672005_4.7uF
*******
.subckt 860160672006_5.6uF 1 2
Rser 1 3 1.36652967282
Lser 2 4 3.637920602E-09
C1 3 4 0.0000056
Rpar 3 4 16666666.6666667
.ends 860160672006_5.6uF
*******
.subckt 860160672007_6.8uF 1 2
Rser 1 3 0.92
Lser 2 4 0.0000000068
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 860160672007_6.8uF
*******
.subckt 860160672008_8.2uF 1 2
Rser 1 3 1.76428312948
Lser 2 4 3.750178848E-09
C1 3 4 0.0000082
Rpar 3 4 12195121.9512195
.ends 860160672008_8.2uF
*******
.subckt 860160672009_10uF 1 2
Rser 1 3 1.60400214929
Lser 2 4 3.334030169E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860160672009_10uF
*******
.subckt 860160672010_15uF 1 2
Rser 1 3 1.40420463201
Lser 2 4 3.962928189E-09
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends 860160672010_15uF
*******
.subckt 860160672011_22uF 1 2
Rser 1 3 1.12048790112
Lser 2 4 4.819832653E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860160672011_22uF
*******
.subckt 860160673012_27uF 1 2
Rser 1 3 0.62317454686
Lser 2 4 3.895436289E-09
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 860160673012_27uF
*******
.subckt 860160673013_33uF 1 2
Rser 1 3 0.624087562311
Lser 2 4 4.915039667E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860160673013_33uF
*******
.subckt 860160673014_39uF 1 2
Rser 1 3 0.37
Lser 2 4 0.0000000072
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860160673014_39uF
*******
.subckt 860160673015_47uF 1 2
Rser 1 3 0.343595281581
Lser 2 4 4.870329504E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860160673015_47uF
*******
.subckt 860160673019_82uF 1 2
Rser 1 3 0.382923990226
Lser 2 4 4.317749582E-09
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860160673019_82uF
*******
.subckt 860160674016_47uF 1 2
Rser 1 3 0.432730094602
Lser 2 4 4.562302287E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860160674016_47uF
*******
.subckt 860160674017_56uF 1 2
Rser 1 3 0.255
Lser 2 4 0.000000008
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860160674017_56uF
*******
.subckt 860160674018_68uF 1 2
Rser 1 3 0.336214692876
Lser 2 4 4.252556875E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860160674018_68uF
*******
.subckt 860160674020_82uF 1 2
Rser 1 3 0.235
Lser 2 4 0.0000000076
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860160674020_82uF
*******
.subckt 860160674021_100uF 1 2
Rser 1 3 0.351996396526
Lser 2 4 4.349817028E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860160674021_100uF
*******
.subckt 860160674022_120uF 1 2
Rser 1 3 0.17
Lser 2 4 0.0000000033
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860160674022_120uF
*******
.subckt 860160674023_150uF 1 2
Rser 1 3 0.145
Lser 2 4 0.000000004
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860160674023_150uF
*******
.subckt 860160674024_180uF 1 2
Rser 1 3 0.118
Lser 2 4 0.0000000032
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160674024_180uF
*******
.subckt 860160675025_180uF 1 2
Rser 1 3 0.183556476718
Lser 2 4 4.577884286E-09
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860160675025_180uF
*******
.subckt 860160675026_220uF 1 2
Rser 1 3 0.111577052239
Lser 2 4 5.430270567E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860160675026_220uF
*******
.subckt 860160675027_270uF 1 2
Rser 1 3 0.10263
Lser 2 4 1.1230117724E-08
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860160675027_270uF
*******
.subckt 860160675028_330uF 1 2
Rser 1 3 0.084
Lser 2 4 0.0000000043
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160675028_330uF
*******
.subckt 860160678029_330uF 1 2
Rser 1 3 0.0692358549308
Lser 2 4 7.788105877E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860160678029_330uF
*******
.subckt 860160678030_470uF 1 2
Rser 1 3 0.057482887837
Lser 2 4 6.977708268E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860160678030_470uF
*******
.subckt 860160678031_560uF 1 2
Rser 1 3 0.0608356632103
Lser 2 4 6.67363026E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860160678031_560uF
*******
.subckt 860160678032_680uF 1 2
Rser 1 3 0.0484110140219
Lser 2 4 8.507066097E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860160678032_680uF
*******
.subckt 860160678033_820uF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000076
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860160678033_820uF
*******
.subckt 860160680034_1mF 1 2
Rser 1 3 0.0382180166321
Lser 2 4 1.3537404135E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 860160680034_1mF
*******
.subckt 860160680035_1.2mF 1 2
Rser 1 3 0.0294035040847
Lser 2 4 1.3334667129E-08
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860160680035_1.2mF
*******
.subckt 860160680036_1.5mF 1 2
Rser 1 3 0.0245785267091
Lser 2 4 1.3296573781E-08
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860160680036_1.5mF
*******
