**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Flat Wire High Current Inductor
* Matchcode:              WE-HCI
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-09
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1030_744323020_0.2u 1 2
Rp 1 2 156.91
Cp 1 2 3.35p
Rs 1 N3 0.00082
L1 N3 2 0.2u
.ends 1030_744323020_0.2u
*******
.subckt 1030_744323033_0.33u 1 2
Rp 1 2 525
Cp 1 2 3.35p
Rs 1 N3 0.00217
L1 N3 2 0.33u
.ends 1030_744323033_0.33u
*******
.subckt 1030_744323056_0.56u 1 2
Rp 1 2 295
Cp 1 2 4.621p
Rs 1 N3 0.00217
L1 N3 2 0.56u
.ends 1030_744323056_0.56u
*******
.subckt 1030_744323068_0.68u 1 2
Rp 1 2 831
Cp 1 2 3.57p
Rs 1 N3 0.00479
L1 N3 2 0.68u
.ends 1030_744323068_0.68u
*******
.subckt 1030_744323100_1u 1 2
Rp 1 2 525
Cp 1 2 4.65p
Rs 1 N3 0.00479
L1 N3 2 1u
.ends 1030_744323100_1u
*******
.subckt 1030_744323120_1.2u 1 2
Rp 1 2 1089
Cp 1 2 5.19p
Rs 1 N3 0.0066
L1 N3 2 1.2u
.ends 1030_744323120_1.2u
*******
.subckt 1030_744323150_1.5u 1 2
Rp 1 2 697
Cp 1 2 6.42p
Rs 1 N3 0.0066
L1 N3 2 1.5u
.ends 1030_744323150_1.5u
*******
.subckt 1030_744323220_2.2u 1 2
Rp 1 2 942
Cp 1 2 5.267p
Rs 1 N3 0.01138
L1 N3 2 2.2u
.ends 1030_744323220_2.2u
*******
.subckt 1040_7443552100_1u 1 2
Rp 1 2 2646
Cp 1 2 3.5p
Rs 1 N3 0.0033
L1 N3 2 1u
.ends 1040_7443552100_1u
*******
.subckt 1040_744355215_0.15u 1 2
Rp 1 2 299.86
Cp 1 2 2.55p
Rs 1 N3 0.00058
L1 N3 2 0.15u
.ends 1040_744355215_0.15u
*******
.subckt 1040_7443552150_1.5u 1 2
Rp 1 2 3213
Cp 1 2 3.63p
Rs 1 N3 0.0053
L1 N3 2 1.5u
.ends 1040_7443552150_1.5u
*******
.subckt 1040_7443552200_2u 1 2
Rp 1 2 605
Cp 1 2 2.59p
Rs 1 N3 0.0073
L1 N3 2 2u
.ends 1040_7443552200_2u
*******
.subckt 1040_7443552280_2.8u 1 2
Rp 1 2 4465
Cp 1 2 4.52p
Rs 1 N3 0.0106
L1 N3 2 2.8u
.ends 1040_7443552280_2.8u
*******
.subckt 1040_744355230_0.3u 1 2
Rp 1 2 1432
Cp 1 2 3.6p
Rs 1 N3 0.0011
L1 N3 2 0.3u
.ends 1040_744355230_0.3u
*******
.subckt 1040_7443552430_4.3u 1 2
Rp 1 2 900
Cp 1 2 3.76p
Rs 1 N3 0.0141
L1 N3 2 4.3u
.ends 1040_7443552430_4.3u
*******
.subckt 1040_744355256_0.56u 1 2
Rp 1 2 2027
Cp 1 2 3.07p
Rs 1 N3 0.00161
L1 N3 2 0.56u
.ends 1040_744355256_0.56u
*******
.subckt 1040_7443552560_5.6u 1 2
Rp 1 2 2725
Cp 1 2 5.3p
Rs 1 N3 0.0206
L1 N3 2 5.6u
.ends 1040_7443552560_5.6u
*******
.subckt 1050_744325016_0.16u 1 2
Rp 1 2 229
Cp 1 2 1.75p
Rs 1 N3 0.00051
L1 N3 2 0.16u
.ends 1050_744325016_0.16u
*******
.subckt 1050_744325040_0.4u 1 2
Rp 1 2 291
Cp 1 2 3.19p
Rs 1 N3 0.00067
L1 N3 2 0.4u
.ends 1050_744325040_0.4u
*******
.subckt 1050_744325072_0.72u 1 2
Rp 1 2 535
Cp 1 2 3.07p
Rs 1 N3 0.0013
L1 N3 2 0.72u
.ends 1050_744325072_0.72u
*******
.subckt 1050_7443251000_10u 1 2
Rp 1 2 2395
Cp 1 2 5.987p
Rs 1 N3 0.0163
L1 N3 2 10u
.ends 1050_7443251000_10u
*******
.subckt 1050_744325120_1.2u 1 2
Rp 1 2 660
Cp 1 2 4.29p
Rs 1 N3 0.0018
L1 N3 2 1.2u
.ends 1050_744325120_1.2u
*******
.subckt 1050_7443251600_16u 1 2
Rp 1 2 4256
Cp 1 2 5.33p
Rs 1 N3 0.0345
L1 N3 2 16u
.ends 1050_7443251600_16u
*******
.subckt 1050_744325180_1.8u 1 2
Rp 1 2 1246
Cp 1 2 3.2p
Rs 1 N3 0.0035
L1 N3 2 1.8u
.ends 1050_744325180_1.8u
*******
.subckt 1050_744325240_2.4u 1 2
Rp 1 2 1099
Cp 1 2 3.83p
Rs 1 N3 0.00475
L1 N3 2 2.4u
.ends 1050_744325240_2.4u
*******
.subckt 1050_744325330_3.3u 1 2
Rp 1 2 1417
Cp 1 2 4.12p
Rs 1 N3 0.0059
L1 N3 2 3.3u
.ends 1050_744325330_3.3u
*******
.subckt 1050_744325420_4.2u 1 2
Rp 1 2 1510
Cp 1 2 4.91p
Rs 1 N3 0.0071
L1 N3 2 4.2u
.ends 1050_744325420_4.2u
*******
.subckt 1050_744325550_5.5u 1 2
Rp 1 2 2100
Cp 1 2 3.89p
Rs 1 N3 0.0103
L1 N3 2 5.5u
.ends 1050_744325550_5.5u
*******
.subckt 1050_744325650_6.5u 1 2
Rp 1 2 1693
Cp 1 2 5.83p
Rs 1 N3 0.0125
L1 N3 2 6.5u
.ends 1050_744325650_6.5u
*******
.subckt 1050_744325780_7.8u 1 2
Rp 1 2 2112
Cp 1 2 6.34p
Rs 1 N3 0.0136
L1 N3 2 7.8u
.ends 1050_744325780_7.8u
*******
.subckt 1335_744313025_0.25u 1 2
Rp 1 2 200
Cp 1 2 3.35p
Rs 1 N3 0.0006
L1 N3 2 0.25u
.ends 1335_744313025_0.25u
*******
.subckt 1335_744313068_0.68u 1 2
Rp 1 2 400
Cp 1 2 5.8p
Rs 1 N3 0.00158
L1 N3 2 0.68u
.ends 1335_744313068_0.68u
*******
.subckt 1335_744313120_1.2u 1 2
Rp 1 2 690
Cp 1 2 6.63p
Rs 1 N3 0.00285
L1 N3 2 1.2u
.ends 1335_744313120_1.2u
*******
.subckt 1335_744313180_1.8u 1 2
Rp 1 2 1079
Cp 1 2 5.35p
Rs 1 N3 0.0056
L1 N3 2 1.8u
.ends 1335_744313180_1.8u
*******
.subckt 1335_744313220_2.2u 1 2
Rp 1 2 914
Cp 1 2 5.75p
Rs 1 N3 0.0057
L1 N3 2 2.2u
.ends 1335_744313220_2.2u
*******
.subckt 1335_744313330_3.3u 1 2
Rp 1 2 1182
Cp 1 2 6p
Rs 1 N3 0.0081
L1 N3 2 3.3u
.ends 1335_744313330_3.3u
*******
.subckt 1350_7443550101_10u 1 2
Rp 1 2 2285
Cp 1 2 9.3p
Rs 1 N3 0.0141
L1 N3 2 10u
.ends 1350_7443550101_10u
*******
.subckt 1350_7443550140_1.4u 1 2
Rp 1 2 1995
Cp 1 2 5.58p
Rs 1 N3 0.0024
L1 N3 2 1.4u
.ends 1350_7443550140_1.4u
*******
.subckt 1350_744355019_0.19u 1 2
Rp 1 2 404
Cp 1 2 1.625p
Rs 1 N3 0.0005
L1 N3 2 0.19u
.ends 1350_744355019_0.19u
*******
.subckt 1350_7443550230_2.3u 1 2
Rp 1 2 2323
Cp 1 2 6p
Rs 1 N3 0.0036
L1 N3 2 2.3u
.ends 1350_7443550230_2.3u
*******
.subckt 1350_7443550320_3.2u 1 2
Rp 1 2 3155
Cp 1 2 5.45p
Rs 1 N3 0.0053
L1 N3 2 3.2u
.ends 1350_7443550320_3.2u
*******
.subckt 1350_744355047_0.47u 1 2
Rp 1 2 720
Cp 1 2 3.56p
Rs 1 N3 0.0009
L1 N3 2 0.47u
.ends 1350_744355047_0.47u
*******
.subckt 1350_7443550480_4.8u 1 2
Rp 1 2 5160
Cp 1 2 4.9p
Rs 1 N3 0.0106
L1 N3 2 4.8u
.ends 1350_7443550480_4.8u
*******
.subckt 1350_7443550600_6u 1 2
Rp 1 2 6000
Cp 1 2 5.3p
Rs 1 N3 0.0137
L1 N3 2 6u
.ends 1350_7443550600_6u
*******
.subckt 1350_7443550820_8.2u 1 2
Rp 1 2 1333
Cp 1 2 9.22p
Rs 1 N3 0.0116
L1 N3 2 8.2u
.ends 1350_7443550820_8.2u
*******
.subckt 1350_744355090_0.9u 1 2
Rp 1 2 1140
Cp 1 2 4.24p
Rs 1 N3 0.00162
L1 N3 2 0.9u
.ends 1350_744355090_0.9u
*******
.subckt 1365_7443551111_11.3u 1 2
Rp 1 2 2457
Cp 1 2 8.47p
Rs 1 N3 0.0091
L1 N3 2 11.3u
.ends 1365_7443551111_11.3u
*******
.subckt 1365_7443551130_1.3u 1 2
Rp 1 2 1750
Cp 1 2 4.4p
Rs 1 N3 0.0017
L1 N3 2 1.3u
.ends 1365_7443551130_1.3u
*******
.subckt 1365_7443551131_13u 1 2
Rp 1 2 2332
Cp 1 2 9.9p
Rs 1 N3 0.011
L1 N3 2 13u
.ends 1365_7443551131_13u
*******
.subckt 1365_7443551151_15.4u 1 2
Rp 1 2 3411
Cp 1 2 8.1p
Rs 1 N3 0.014
L1 N3 2 15.4u
.ends 1365_7443551151_15.4u
*******
.subckt 1365_7443551181_18u 1 2
Rp 1 2 5179
Cp 1 2 5.65p
Rs 1 N3 0.022
L1 N3 2 18u
.ends 1365_7443551181_18u
*******
.subckt 1365_7443551200_2u 1 2
Rp 1 2 2270
Cp 1 2 4.9p
Rs 1 N3 0.0025
L1 N3 2 2u
.ends 1365_7443551200_2u
*******
.subckt 1365_744355122_0.2u 1 2
Rp 1 2 400
Cp 1 2 1.67p
Rs 1 N3 0.00037
L1 N3 2 0.2u
.ends 1365_744355122_0.2u
*******
.subckt 1365_7443551221_22u 1 2
Rp 1 2 4310
Cp 1 2 6.2p
Rs 1 N3 0.0247
L1 N3 2 22u
.ends 1365_7443551221_22u
*******
.subckt 1365_7443551280_2.8u 1 2
Rp 1 2 3044
Cp 1 2 5.1p
Rs 1 N3 0.0034
L1 N3 2 2.8u
.ends 1365_7443551280_2.8u
*******
.subckt 1365_7443551331_33u 1 2
Rp 1 2 5276
Cp 1 2 7.71p
Rs 1 N3 0.0305
L1 N3 2 33u
.ends 1365_7443551331_33u
*******
.subckt 1365_7443551370_3.7u 1 2
Rp 1 2 3948
Cp 1 2 5.02p
Rs 1 N3 0.0049
L1 N3 2 3.7u
.ends 1365_7443551370_3.7u
*******
.subckt 1365_744355147_0.47u 1 2
Rp 1 2 706
Cp 1 2 4p
Rs 1 N3 0.00064
L1 N3 2 0.47u
.ends 1365_744355147_0.47u
*******
.subckt 1365_7443551470_4.7u 1 2
Rp 1 2 5393
Cp 1 2 4.4p
Rs 1 N3 0.0069
L1 N3 2 4.7u
.ends 1365_7443551470_4.7u
*******
.subckt 1365_7443551600_6u 1 2
Rp 1 2 6676
Cp 1 2 4.1p
Rs 1 N3 0.0083
L1 N3 2 6u
.ends 1365_7443551600_6u
*******
.subckt 1365_7443551730_7.3u 1 2
Rp 1 2 2435
Cp 1 2 5.45p
Rs 1 N3 0.0059
L1 N3 2 7.3u
.ends 1365_7443551730_7.3u
*******
.subckt 1365_744355182_0.82u 1 2
Rp 1 2 1173
Cp 1 2 5.38p
Rs 1 N3 0.00104
L1 N3 2 0.82u
.ends 1365_744355182_0.82u
*******
.subckt 1365_7443551920_9.2u 1 2
Rp 1 2 2657
Cp 1 2 6.6p
Rs 1 N3 0.0076
L1 N3 2 9.2u
.ends 1365_7443551920_9.2u
*******
.subckt 1890_7443556082_0.82u 1 2
Rp 1 2 270
Cp 1 2 6.35p
Rs 1 N3 0.00054
L1 N3 2 0.82u
.ends 1890_7443556082_0.82u
*******
.subckt 1890_74435561100_10u 1 2
Rp 1 2 1459
Cp 1 2 9.409p
Rs 1 N3 0.0069
L1 N3 2 10u
.ends 1890_74435561100_10u
*******
.subckt 1890_7443556130_1.3u 1 2
Rp 1 2 349
Cp 1 2 6.13p
Rs 1 N3 0.00094
L1 N3 2 1.3u
.ends 1890_7443556130_1.3u
*******
.subckt 1890_7443556190_1.9u 1 2
Rp 1 2 464
Cp 1 2 6.816p
Rs 1 N3 0.0012
L1 N3 2 1.9u
.ends 1890_7443556190_1.9u
*******
.subckt 1890_7443556260_2.6u 1 2
Rp 1 2 626
Cp 1 2 6.508p
Rs 1 N3 0.00158
L1 N3 2 2.6u
.ends 1890_7443556260_2.6u
*******
.subckt 1890_7443556350_3.5u 1 2
Rp 1 2 735
Cp 1 2 6.17p
Rs 1 N3 0.0031
L1 N3 2 3.5u
.ends 1890_7443556350_3.5u
*******
.subckt 1890_7443556450_4.5u 1 2
Rp 1 2 1050
Cp 1 2 6.45p
Rs 1 N3 0.0034
L1 N3 2 4.5u
.ends 1890_7443556450_4.5u
*******
.subckt 1890_7443556560_5.6u 1 2
Rp 1 2 1071
Cp 1 2 7.138p
Rs 1 N3 0.0037
L1 N3 2 5.6u
.ends 1890_7443556560_5.6u
*******
.subckt 1890_7443556680_6.8u 1 2
Rp 1 2 1186
Cp 1 2 8.508p
Rs 1 N3 0.0041
L1 N3 2 6.8u
.ends 1890_7443556680_6.8u
*******
.subckt 1890_74435571100_10u 1 2
Rp 1 2 2300
Cp 1 2 14p
Rs 1 N3 0.0069
L1 N3 2 10u
.ends 1890_74435571100_10u
*******
.subckt 1890_74435571500_15u 1 2
Rp 1 2 2340
Cp 1 2 16.87p
Rs 1 N3 0.009
L1 N3 2 15u
.ends 1890_74435571500_15u
*******
.subckt 1890_74435572200_22u 1 2
Rp 1 2 4220
Cp 1 2 14.91p
Rs 1 N3 0.0146
L1 N3 2 22u
.ends 1890_74435572200_22u
*******
.subckt 1890_74435573300_33u 1 2
Rp 1 2 4860
Cp 1 2 11.6p
Rs 1 N3 0.0217
L1 N3 2 33u
.ends 1890_74435573300_33u
*******
.subckt 1890_74435574700_47u 1 2
Rp 1 2 13200
Cp 1 2 17.78p
Rs 1 N3 0.0335
L1 N3 2 47u
.ends 1890_74435574700_47u
*******
.subckt 1890_7443557560_5.6u 1 2
Rp 1 2 1671
Cp 1 2 9.043p
Rs 1 N3 0.00274
L1 N3 2 5.6u
.ends 1890_7443557560_5.6u
*******
.subckt 1890_7443557760_7.6u 1 2
Rp 1 2 1980
Cp 1 2 9.893p
Rs 1 N3 0.0037
L1 N3 2 7.6u
.ends 1890_7443557760_7.6u
*******
.subckt 2212_74435580330_3.3u 1 2
Rp 1 2 1831
Cp 1 2 8.401p
Rs 1 N3 0.0017
L1 N3 2 3.3u
.ends 2212_74435580330_3.3u
*******
.subckt 5040_744316022_0.22u 1 2
Rp 1 2 190.171
Cp 1 2 1.527p
Rs 1 N3 0.00125
L1 N3 2 0.22u
.ends 5040_744316022_0.22u
*******
.subckt 5040_744316033_0.33u 1 2
Rp 1 2 191.468
Cp 1 2 1.36p
Rs 1 N3 0.00175
L1 N3 2 0.33u
.ends 5040_744316033_0.33u
*******
.subckt 5040_744316047_0.47u 1 2
Rp 1 2 276.518
Cp 1 2 1.652p
Rs 1 N3 0.00275
L1 N3 2 0.47u
.ends 5040_744316047_0.47u
*******
.subckt 5040_744316068_0.68u 1 2
Rp 1 2 395.249
Cp 1 2 1.382p
Rs 1 N3 0.004
L1 N3 2 0.68u
.ends 5040_744316068_0.68u
*******
.subckt 5040_744316100_1u 1 2
Rp 1 2 530.165
Cp 1 2 2.021p
Rs 1 N3 0.00475
L1 N3 2 1u
.ends 5040_744316100_1u
*******
.subckt 5040_744316150_1.5u 1 2
Rp 1 2 692.752
Cp 1 2 2.226p
Rs 1 N3 0.00815
L1 N3 2 1.5u
.ends 5040_744316150_1.5u
*******
.subckt 5040_744316220_2.2u 1 2
Rp 1 2 846.631
Cp 1 2 1.821p
Rs 1 N3 0.0113
L1 N3 2 2.2u
.ends 5040_744316220_2.2u
*******
.subckt 5040_744316330_3.3u 1 2
Rp 1 2 1519.2
Cp 1 2 2.413p
Rs 1 N3 0.0185
L1 N3 2 3.3u
.ends 5040_744316330_3.3u
*******
.subckt 5040_744316470_4.7u 1 2
Rp 1 2 1365.6
Cp 1 2 2.51p
Rs 1 N3 0.0245
L1 N3 2 4.7u
.ends 5040_744316470_4.7u
*******
.subckt 5040_744316560_5.6u 1 2
Rp 1 2 1377.89
Cp 1 2 3.087p
Rs 1 N3 0.0285
L1 N3 2 5.6u
.ends 5040_744316560_5.6u
*******
.subckt 7030_744310013_0.13u 1 2
Rp 1 2 207
Cp 1 2 0.68p
Rs 1 N3 0.00091
L1 N3 2 0.13u
.ends 7030_744310013_0.13u
*******
.subckt 7030_744310024_0.24u 1 2
Rp 1 2 368
Cp 1 2 1.05p
Rs 1 N3 0.0018
L1 N3 2 0.24u
.ends 7030_744310024_0.24u
*******
.subckt 7030_744310055_0.52u 1 2
Rp 1 2 500
Cp 1 2 1.25p
Rs 1 N3 0.0037
L1 N3 2 0.52u
.ends 7030_744310055_0.52u
*******
.subckt 7030_744310095_0.95u 1 2
Rp 1 2 720
Cp 1 2 1.17p
Rs 1 N3 0.0062
L1 N3 2 0.95u
.ends 7030_744310095_0.95u
*******
.subckt 7030_744310115_1.15u 1 2
Rp 1 2 933
Cp 1 2 1.24p
Rs 1 N3 0.0086
L1 N3 2 1.15u
.ends 7030_744310115_1.15u
*******
.subckt 7030_744310150_1.5u 1 2
Rp 1 2 695
Cp 1 2 2.72p
Rs 1 N3 0.0127
L1 N3 2 1.5u
.ends 7030_744310150_1.5u
*******
.subckt 7030_744310200_2u 1 2
Rp 1 2 1120
Cp 1 2 1.6p
Rs 1 N3 0.0142
L1 N3 2 2u
.ends 7030_744310200_2u
*******
.subckt 7040_744311022_0.22u 1 2
Rp 1 2 262
Cp 1 2 2p
Rs 1 N3 0.0011
L1 N3 2 0.22u
.ends 7040_744311022_0.22u
*******
.subckt 7040_744311047_0.4u 1 2
Rp 1 2 506
Cp 1 2 1.57p
Rs 1 N3 0.00185
L1 N3 2 0.4u
.ends 7040_744311047_0.4u
*******
.subckt 7040_744311068_0.68u 1 2
Rp 1 2 732
Cp 1 2 1.02p
Rs 1 N3 0.0031
L1 N3 2 0.68u
.ends 7040_744311068_0.68u
*******
.subckt 7040_744311100_1u 1 2
Rp 1 2 756
Cp 1 2 2.85p
Rs 1 N3 0.0046
L1 N3 2 1u
.ends 7040_744311100_1u
*******
.subckt 7040_744311150_1.5u 1 2
Rp 1 2 1212
Cp 1 2 1.18p
Rs 1 N3 0.0066
L1 N3 2 1.5u
.ends 7040_744311150_1.5u
*******
.subckt 7040_744311220_2.2u 1 2
Rp 1 2 1495
Cp 1 2 1.19p
Rs 1 N3 0.0114
L1 N3 2 2.2u
.ends 7040_744311220_2.2u
*******
.subckt 7040_744311330_3.3u 1 2
Rp 1 2 2464
Cp 1 2 1.81p
Rs 1 N3 0.0172
L1 N3 2 3.3u
.ends 7040_744311330_3.3u
*******
.subckt 7040_744311470_4.7u 1 2
Rp 1 2 2575
Cp 1 2 1.81p
Rs 1 N3 0.0195
L1 N3 2 4.7u
.ends 7040_744311470_4.7u
*******
.subckt 7050_744314024_0.24u 1 2
Rp 1 2 220
Cp 1 2 1.95p
Rs 1 N3 0.001
L1 N3 2 0.24u
.ends 7050_744314024_0.24u
*******
.subckt 7050_744314047_0.47u 1 2
Rp 1 2 372
Cp 1 2 1.78p
Rs 1 N3 0.00135
L1 N3 2 0.47u
.ends 7050_744314047_0.47u
*******
.subckt 7050_744314076_0.76u 1 2
Rp 1 2 588
Cp 1 2 1.62p
Rs 1 N3 0.00225
L1 N3 2 0.76u
.ends 7050_744314076_0.76u
*******
.subckt 7050_744314101_10u 1 2
Rp 1 2 3803
Cp 1 2 2.03p
Rs 1 N3 0.033
L1 N3 2 10u
.ends 7050_744314101_10u
*******
.subckt 7050_744314110_1.1u 1 2
Rp 1 2 810
Cp 1 2 1.61p
Rs 1 N3 0.00315
L1 N3 2 1.1u
.ends 7050_744314110_1.1u
*******
.subckt 7050_744314150_1.5u 1 2
Rp 1 2 820
Cp 1 2 2.11p
Rs 1 N3 0.0043
L1 N3 2 1.5u
.ends 7050_744314150_1.5u
*******
.subckt 7050_744314200_2u 1 2
Rp 1 2 1356
Cp 1 2 3.37p
Rs 1 N3 0.00585
L1 N3 2 2u
.ends 7050_744314200_2u
*******
.subckt 7050_744314330_3.3u 1 2
Rp 1 2 1694
Cp 1 2 2.18p
Rs 1 N3 0.009
L1 N3 2 3.3u
.ends 7050_744314330_3.3u
*******
.subckt 7050_744314490_4.9u 1 2
Rp 1 2 1732
Cp 1 2 2.15p
Rs 1 N3 0.0145
L1 N3 2 4.9u
.ends 7050_744314490_4.9u
*******
.subckt 7050_744314650_6.5u 1 2
Rp 1 2 2330
Cp 1 2 2p
Rs 1 N3 0.0215
L1 N3 2 6.5u
.ends 7050_744314650_6.5u
*******
.subckt 7050_744314760_7.6u 1 2
Rp 1 2 3119
Cp 1 2 2.03p
Rs 1 N3 0.0302
L1 N3 2 7.6u
.ends 7050_744314760_7.6u
*******
.subckt 7050_744314850_8.5u 1 2
Rp 1 2 3563
Cp 1 2 1.9p
Rs 1 N3 0.0325
L1 N3 2 8.5u
.ends 7050_744314850_8.5u
*******
.subckt 2212_74435580680_6.8u 1 2
Rp 1 2 1900
Cp 1 2 9.78p
Rs 1 N3 0.0021
L1 N3 2 6.8u
.ends 2212_74435580680_6.8u
*******
.subckt 2212_74435580820_8.2u 1 2
Rp 1 2 2350
Cp 1 2 10p
Rs 1 N3 0.0027
L1 N3 2 8.2u
.ends 2212_74435580820_8.2u
*******
.subckt 2212_74435581000_10u 1 2
Rp 1 2 2833
Cp 1 2 9p
Rs 1 N3 0.0034
L1 N3 2 10u
.ends 2212_74435581000_10u
*******
.subckt 2212_74435581200_12u 1 2
Rp 1 2 3150
Cp 1 2 9.5p
Rs 1 N3 0.0043
L1 N3 2 12u
.ends 2212_74435581200_12u
*******
.subckt 2212_74435582200_22u 1 2
Rp 1 2 3500
Cp 1 2 16p
Rs 1 N3 0.007
L1 N3 2 22u
.ends 2212_74435582200_22u
*******
.subckt 2212_74435583300_33u 1 2
Rp 1 2 7500
Cp 1 2 11p
Rs 1 N3 0.0132
L1 N3 2 33u
.ends 2212_74435583300_33u
*******
.subckt 2212_74435584700_47u 1 2
Rp 1 2 9000
Cp 1 2 13p
Rs 1 N3 0.0192
L1 N3 2 47u
.ends 2212_74435584700_47u
*******
.subckt 2212_74435586800_68u 1 2
Rp 1 2 12000
Cp 1 2 11p
Rs 1 N3 0.0273
L1 N3 2 68u
.ends 2212_74435586800_68u
*******
.subckt 2212_74435588200_82u 1 2
Rp 1 2 13250
Cp 1 2 12p
Rs 1 N3 0.0304
L1 N3 2 82u
.ends 2212_74435588200_82u
*******
