**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Tiny Power Inductor
* Matchcode:              WE-TPC 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1028_744065001_1u 1 2
Rp 1 2 1445
Cp 1 2 2.32p
Rs 1 N3 0.0049
L1 N3 2 1u
.ends 1028_744065001_1u
*******
.subckt 1028_7440650015_1.5u 1 2
Rp 1 2 2272
Cp 1 2 2.24p
Rs 1 N3 0.0073
L1 N3 2 1.5u
.ends 1028_7440650015_1.5u
*******
.subckt 1028_7440650022_2.2u 1 2
Rp 1 2 3170
Cp 1 2 2.46p
Rs 1 N3 0.011
L1 N3 2 2.2u
.ends 1028_7440650022_2.2u
*******
.subckt 1028_7440650033_3.3u 1 2
Rp 1 2 3402
Cp 1 2 2.53p
Rs 1 N3 0.015
L1 N3 2 3.3u
.ends 1028_7440650033_3.3u
*******
.subckt 1028_7440650047_4.7u 1 2
Rp 1 2 5922
Cp 1 2 2.74p
Rs 1 N3 0.0165
L1 N3 2 4.7u
.ends 1028_7440650047_4.7u
*******
.subckt 1028_7440650068_6.8u 1 2
Rp 1 2 6495
Cp 1 2 2.95p
Rs 1 N3 0.025
L1 N3 2 6.8u
.ends 1028_7440650068_6.8u
*******
.subckt 1028_7440650082_8.2u 1 2
Rp 1 2 8057
Cp 1 2 2.79p
Rs 1 N3 0.0285
L1 N3 2 8.2u
.ends 1028_7440650082_8.2u
*******
.subckt 1028_744065100_10u 1 2
Rp 1 2 9830
Cp 1 2 2.92p
Rs 1 N3 0.04
L1 N3 2 10u
.ends 1028_744065100_10u
*******
.subckt 1028_744065101_100u 1 2
Rp 1 2 49583
Cp 1 2 2.82p
Rs 1 N3 0.365
L1 N3 2 100u
.ends 1028_744065101_100u
*******
.subckt 1028_744065121_120u 1 2
Rp 1 2 54931
Cp 1 2 3.38p
Rs 1 N3 0.428
L1 N3 2 120u
.ends 1028_744065121_120u
*******
.subckt 1028_744065150_15u 1 2
Rp 1 2 12382
Cp 1 2 2.36p
Rs 1 N3 0.069
L1 N3 2 15u
.ends 1028_744065150_15u
*******
.subckt 1028_744065151_150u 1 2
Rp 1 2 49255
Cp 1 2 3.7p
Rs 1 N3 0.53
L1 N3 2 150u
.ends 1028_744065151_150u
*******
.subckt 1028_744065220_22u 1 2
Rp 1 2 15135
Cp 1 2 3.48p
Rs 1 N3 0.104
L1 N3 2 22u
.ends 1028_744065220_22u
*******
.subckt 1028_744065221_220u 1 2
Rp 1 2 56966
Cp 1 2 3.738p
Rs 1 N3 0.75
L1 N3 2 220u
.ends 1028_744065221_220u
*******
.subckt 1028_744065330_33u 1 2
Rp 1 2 21315
Cp 1 2 2.7p
Rs 1 N3 0.139
L1 N3 2 33u
.ends 1028_744065330_33u
*******
.subckt 1028_744065470_47u 1 2
Rp 1 2 26383
Cp 1 2 2.86p
Rs 1 N3 0.167
L1 N3 2 47u
.ends 1028_744065470_47u
*******
.subckt 1028_744065560_56u 1 2
Rp 1 2 28460
Cp 1 2 3.12p
Rs 1 N3 0.208
L1 N3 2 56u
.ends 1028_744065560_56u
*******
.subckt 1028_744065680_68u 1 2
Rp 1 2 32141
Cp 1 2 3.41p
Rs 1 N3 0.232
L1 N3 2 68u
.ends 1028_744065680_68u
*******
.subckt 1028_744065820_82u 1 2
Rp 1 2 44443
Cp 1 2 3.2p
Rs 1 N3 0.323
L1 N3 2 82u
.ends 1028_744065820_82u
*******
.subckt 1038_7440660015_1.5u 1 2
Rp 1 2 2495
Cp 1 2 3.57p
Rs 1 N3 0.0052
L1 N3 2 1.5u
.ends 1038_7440660015_1.5u
*******
.subckt 1038_7440660022_2.2u 1 2
Rp 1 2 3200
Cp 1 2 3.2p
Rs 1 N3 0.0077
L1 N3 2 2.2u
.ends 1038_7440660022_2.2u
*******
.subckt 1038_7440660035_3.5u 1 2
Rp 1 2 5448
Cp 1 2 3.9p
Rs 1 N3 0.0115
L1 N3 2 3.5u
.ends 1038_7440660035_3.5u
*******
.subckt 1038_744066005_5u 1 2
Rp 1 2 5450
Cp 1 2 3.3p
Rs 1 N3 0.0145
L1 N3 2 5u
.ends 1038_744066005_5u
*******
.subckt 1038_7440660062_6.2u 1 2
Rp 1 2 6602
Cp 1 2 4.52p
Rs 1 N3 0.0165
L1 N3 2 6.2u
.ends 1038_7440660062_6.2u
*******
.subckt 1038_744066100_10u 1 2
Rp 1 2 8190
Cp 1 2 4.17p
Rs 1 N3 0.025
L1 N3 2 10u
.ends 1038_744066100_10u
*******
.subckt 1038_744066101_100u 1 2
Rp 1 2 45371
Cp 1 2 5p
Rs 1 N3 0.255
L1 N3 2 100u
.ends 1038_744066101_100u
*******
.subckt 1038_744066150_15u 1 2
Rp 1 2 11832
Cp 1 2 4.13p
Rs 1 N3 0.037
L1 N3 2 15u
.ends 1038_744066150_15u
*******
.subckt 1038_744066151_150u 1 2
Rp 1 2 53241
Cp 1 2 4.95p
Rs 1 N3 0.35
L1 N3 2 150u
.ends 1038_744066151_150u
*******
.subckt 1038_744066180_18u 1 2
Rp 1 2 14535
Cp 1 2 4.94p
Rs 1 N3 0.054
L1 N3 2 18u
.ends 1038_744066180_18u
*******
.subckt 1038_744066220_22u 1 2
Rp 1 2 12878
Cp 1 2 5.36p
Rs 1 N3 0.0558
L1 N3 2 22u
.ends 1038_744066220_22u
*******
.subckt 1038_744066221_220u 1 2
Rp 1 2 58000
Cp 1 2 5p
Rs 1 N3 0.57
L1 N3 2 220u
.ends 1038_744066221_220u
*******
.subckt 1038_744066330_33u 1 2
Rp 1 2 20600
Cp 1 2 4.58p
Rs 1 N3 0.092
L1 N3 2 33u
.ends 1038_744066330_33u
*******
.subckt 1038_744066331_330u 1 2
Rp 1 2 107820
Cp 1 2 5.45p
Rs 1 N3 0.77
L1 N3 2 330u
.ends 1038_744066331_330u
*******
.subckt 1038_744066470_47u 1 2
Rp 1 2 25640
Cp 1 2 6.17p
Rs 1 N3 0.121
L1 N3 2 47u
.ends 1038_744066470_47u
*******
.subckt 1038_744066680_68u 1 2
Rp 1 2 33120
Cp 1 2 5.7p
Rs 1 N3 0.185
L1 N3 2 68u
.ends 1038_744066680_68u
*******
.subckt 1038_744066681_680u 1 2
Rp 1 2 116034
Cp 1 2 6.25p
Rs 1 N3 1.65
L1 N3 2 680u
.ends 1038_744066681_680u
*******
.subckt 2811_744028000056_0.056u 1 2
Rp 1 2 123
Cp 1 2 0.03p
Rs 1 N3 0.0115
L1 N3 2 0.056u
.ends 2811_744028000056_0.056u
*******
.subckt 2811_74402800015_0.15u 1 2
Rp 1 2 290
Cp 1 2 0.19p
Rs 1 N3 0.018
L1 N3 2 0.15u
.ends 2811_74402800015_0.15u
*******
.subckt 2811_74402800033_0.33u 1 2
Rp 1 2 578
Cp 1 2 0.265p
Rs 1 N3 0.027
L1 N3 2 0.33u
.ends 2811_74402800033_0.33u
*******
.subckt 2811_74402800047_0.47u 1 2
Rp 1 2 883
Cp 1 2 0.432p
Rs 1 N3 0.036
L1 N3 2 0.47u
.ends 2811_74402800047_0.47u
*******
.subckt 2811_74402800082_0.82u 1 2
Rp 1 2 1833
Cp 1 2 0.512p
Rs 1 N3 0.053
L1 N3 2 0.82u
.ends 2811_74402800082_0.82u
*******
.subckt 2811_744028001_1u 1 2
Rp 1 2 2000
Cp 1 2 1.55p
Rs 1 N3 0.065
L1 N3 2 1u
.ends 2811_744028001_1u
*******
.subckt 2811_744028002_2.2u 1 2
Rp 1 2 2900
Cp 1 2 1.77p
Rs 1 N3 0.125
L1 N3 2 2.2u
.ends 2811_744028002_2.2u
*******
.subckt 2811_744028003_3.3u 1 2
Rp 1 2 5210
Cp 1 2 1.53p
Rs 1 N3 0.185
L1 N3 2 3.3u
.ends 2811_744028003_3.3u
*******
.subckt 2811_744028004_4.7u 1 2
Rp 1 2 5570
Cp 1 2 1.69p
Rs 1 N3 0.265
L1 N3 2 4.7u
.ends 2811_744028004_4.7u
*******
.subckt 2811_744028006_6.8u 1 2
Rp 1 2 6760
Cp 1 2 1.54p
Rs 1 N3 0.325
L1 N3 2 6.8u
.ends 2811_744028006_6.8u
*******
.subckt 2813_744029000068_0.068u 1 2
Rp 1 2 260
Cp 1 2 0.03p
Rs 1 N3 0.0105
L1 N3 2 0.068u
.ends 2813_744029000068_0.068u
*******
.subckt 2813_74402900016_0.16u 1 2
Rp 1 2 432
Cp 1 2 0.18p
Rs 1 N3 0.016
L1 N3 2 0.16u
.ends 2813_74402900016_0.16u
*******
.subckt 2813_74402900033_0.33u 1 2
Rp 1 2 533
Cp 1 2 0.254p
Rs 1 N3 0.023
L1 N3 2 0.33u
.ends 2813_74402900033_0.33u
*******
.subckt 2813_74402900047_0.47u 1 2
Rp 1 2 836
Cp 1 2 0.43p
Rs 1 N3 0.029
L1 N3 2 0.47u
.ends 2813_74402900047_0.47u
*******
.subckt 2813_74402900082_0.82u 1 2
Rp 1 2 1632
Cp 1 2 0.541p
Rs 1 N3 0.036
L1 N3 2 0.82u
.ends 2813_74402900082_0.82u
*******
.subckt 2813_744029001_1u 1 2
Rp 1 2 1550
Cp 1 2 1.63p
Rs 1 N3 0.045
L1 N3 2 1u
.ends 2813_744029001_1u
*******
.subckt 2813_744029002_2.2u 1 2
Rp 1 2 3300
Cp 1 2 1.7p
Rs 1 N3 0.088
L1 N3 2 2.2u
.ends 2813_744029002_2.2u
*******
.subckt 2813_744029003_3.3u 1 2
Rp 1 2 3900
Cp 1 2 1.7p
Rs 1 N3 0.11
L1 N3 2 3.3u
.ends 2813_744029003_3.3u
*******
.subckt 2813_744029004_4.7u 1 2
Rp 1 2 6000
Cp 1 2 1.65p
Rs 1 N3 0.17
L1 N3 2 4.7u
.ends 2813_744029004_4.7u
*******
.subckt 2813_744029006_6.8u 1 2
Rp 1 2 5900
Cp 1 2 1.9p
Rs 1 N3 0.25
L1 N3 2 6.8u
.ends 2813_744029006_6.8u
*******
.subckt 2813_744029100_10u 1 2
Rp 1 2 10000
Cp 1 2 1.725p
Rs 1 N3 0.39
L1 N3 2 10u
.ends 2813_744029100_10u
*******
.subckt 2828_74402500030_0.3u 1 2
Rp 1 2 300
Cp 1 2 0.885p
Rs 1 N3 0.015
L1 N3 2 0.3u
.ends 2828_74402500030_0.3u
*******
.subckt 2828_74402500047_0.47u 1 2
Rp 1 2 477
Cp 1 2 0.816p
Rs 1 N3 0.019
L1 N3 2 0.47u
.ends 2828_74402500047_0.47u
*******
.subckt 2828_74402500072_0.72u 1 2
Rp 1 2 600
Cp 1 2 0.966p
Rs 1 N3 0.0235
L1 N3 2 0.72u
.ends 2828_74402500072_0.72u
*******
.subckt 2828_744025001_1.2u 1 2
Rp 1 2 850
Cp 1 2 1.128p
Rs 1 N3 0.036
L1 N3 2 1.2u
.ends 2828_744025001_1.2u
*******
.subckt 2828_744025002_2.2u 1 2
Rp 1 2 1700
Cp 1 2 1.3p
Rs 1 N3 0.057
L1 N3 2 2.2u
.ends 2828_744025002_2.2u
*******
.subckt 2828_744025003_3.3u 1 2
Rp 1 2 2500
Cp 1 2 1.8p
Rs 1 N3 0.085
L1 N3 2 3.3u
.ends 2828_744025003_3.3u
*******
.subckt 2828_744025004_4.7u 1 2
Rp 1 2 3800
Cp 1 2 2.5p
Rs 1 N3 0.1
L1 N3 2 4.7u
.ends 2828_744025004_4.7u
*******
.subckt 2828_744025006_6.8u 1 2
Rp 1 2 3303
Cp 1 2 1.699p
Rs 1 N3 0.142
L1 N3 2 6.8u
.ends 2828_744025006_6.8u
*******
.subckt 2828_744025100_10u 1 2
Rp 1 2 6412
Cp 1 2 2.33p
Rs 1 N3 0.17
L1 N3 2 10u
.ends 2828_744025100_10u
*******
.subckt 2828_744025150_15u 1 2
Rp 1 2 10373
Cp 1 2 1.734p
Rs 1 N3 0.356
L1 N3 2 15u
.ends 2828_744025150_15u
*******
.subckt 2828_744025220_22u 1 2
Rp 1 2 13000
Cp 1 2 2.815p
Rs 1 N3 0.525
L1 N3 2 22u
.ends 2828_744025220_22u
*******
.subckt 2828_744025270_27u 1 2
Rp 1 2 10349
Cp 1 2 4.699p
Rs 1 N3 0.745
L1 N3 2 27u
.ends 2828_744025270_27u
*******
.subckt 2828_744025330_33u 1 2
Rp 1 2 12077
Cp 1 2 6p
Rs 1 N3 0.84
L1 N3 2 33u
.ends 2828_744025330_33u
*******
.subckt 3510_744030001_1.2u 1 2
Rp 1 2 2690
Cp 1 2 0.52p
Rs 1 N3 0.095
L1 N3 2 1.2u
.ends 3510_744030001_1.2u
*******
.subckt 3510_744030002_2.2u 1 2
Rp 1 2 4065
Cp 1 2 0.575p
Rs 1 N3 0.14
L1 N3 2 2.2u
.ends 3510_744030002_2.2u
*******
.subckt 3510_744030003_3.3u 1 2
Rp 1 2 6383
Cp 1 2 0.693p
Rs 1 N3 0.198
L1 N3 2 3.3u
.ends 3510_744030003_3.3u
*******
.subckt 3510_744030004_4.7u 1 2
Rp 1 2 7861
Cp 1 2 0.589p
Rs 1 N3 0.252
L1 N3 2 4.7u
.ends 3510_744030004_4.7u
*******
.subckt 3510_7440300047_0.47u 1 2
Rp 1 2 1110
Cp 1 2 1.739p
Rs 1 N3 0.048
L1 N3 2 0.47u
.ends 3510_7440300047_0.47u
*******
.subckt 3510_744030006_6.8u 1 2
Rp 1 2 9968
Cp 1 2 0.676p
Rs 1 N3 0.4
L1 N3 2 6.8u
.ends 3510_744030006_6.8u
*******
.subckt 3510_7440300068_0.68u 1 2
Rp 1 2 1494
Cp 1 2 1.754p
Rs 1 N3 0.06
L1 N3 2 0.68u
.ends 3510_7440300068_0.68u
*******
.subckt 3816_744031001_1.5u 1 2
Rp 1 2 2272
Cp 1 2 0.974p
Rs 1 N3 0.04
L1 N3 2 1.5u
.ends 3816_744031001_1.5u
*******
.subckt 3816_744031002_2.5u 1 2
Rp 1 2 4428
Cp 1 2 1.15p
Rs 1 N3 0.05
L1 N3 2 2.5u
.ends 3816_744031002_2.5u
*******
.subckt 3816_744031003_3.6u 1 2
Rp 1 2 4823
Cp 1 2 0.944p
Rs 1 N3 0.066
L1 N3 2 3.6u
.ends 3816_744031003_3.6u
*******
.subckt 3816_744031004_4.7u 1 2
Rp 1 2 5904
Cp 1 2 1.235p
Rs 1 N3 0.09
L1 N3 2 4.7u
.ends 3816_744031004_4.7u
*******
.subckt 3816_7440310047_0.47u 1 2
Rp 1 2 574
Cp 1 2 1.727p
Rs 1 N3 0.016
L1 N3 2 0.47u
.ends 3816_7440310047_0.47u
*******
.subckt 3816_744031006_6.8u 1 2
Rp 1 2 6886
Cp 1 2 1.067p
Rs 1 N3 0.135
L1 N3 2 6.8u
.ends 3816_744031006_6.8u
*******
.subckt 3816_744031010_1u 1 2
Rp 1 2 1309
Cp 1 2 2.138p
Rs 1 N3 0.026
L1 N3 2 1u
.ends 3816_744031010_1u
*******
.subckt 3816_744031100_10u 1 2
Rp 1 2 10770
Cp 1 2 1.28p
Rs 1 N3 0.185
L1 N3 2 10u
.ends 3816_744031100_10u
*******
.subckt 3816_744031101_100u 1 2
Rp 1 2 43423
Cp 1 2 1.37p
Rs 1 N3 1.93
L1 N3 2 100u
.ends 3816_744031101_100u
*******
.subckt 3816_744031150_15u 1 2
Rp 1 2 11900
Cp 1 2 1.35p
Rs 1 N3 0.255
L1 N3 2 15u
.ends 3816_744031150_15u
*******
.subckt 3816_744031220_22u 1 2
Rp 1 2 14548
Cp 1 2 1.388p
Rs 1 N3 0.41
L1 N3 2 22u
.ends 3816_744031220_22u
*******
.subckt 3816_744031330_33u 1 2
Rp 1 2 15045
Cp 1 2 2.413p
Rs 1 N3 0.635
L1 N3 2 33u
.ends 3816_744031330_33u
*******
.subckt 3816_744031470_47u 1 2
Rp 1 2 42811
Cp 1 2 1.34p
Rs 1 N3 0.94
L1 N3 2 47u
.ends 3816_744031470_47u
*******
.subckt 3816_744031680_68u 1 2
Rp 1 2 43152
Cp 1 2 1.36p
Rs 1 N3 1.15
L1 N3 2 68u
.ends 3816_744031680_68u
*******
.subckt 4818_74404200056_0.56u 1 2
Rp 1 2 947
Cp 1 2 1.776p
Rs 1 N3 0.019
L1 N3 2 0.56u
.ends 4818_74404200056_0.56u
*******
.subckt 4818_744042001_1u 1 2
Rp 1 2 1444
Cp 1 2 0.518p
Rs 1 N3 0.02
L1 N3 2 1u
.ends 4818_744042001_1u
*******
.subckt 4818_7440420018_1.8u 1 2
Rp 1 2 2627
Cp 1 2 1.322p
Rs 1 N3 0.04
L1 N3 2 1.8u
.ends 4818_7440420018_1.8u
*******
.subckt 4818_7440420027_2.7u 1 2
Rp 1 2 3189
Cp 1 2 1.17p
Rs 1 N3 0.047
L1 N3 2 2.7u
.ends 4818_7440420027_2.7u
*******
.subckt 4818_744042003_3.3u 1 2
Rp 1 2 3960
Cp 1 2 1.227p
Rs 1 N3 0.05
L1 N3 2 3.3u
.ends 4818_744042003_3.3u
*******
.subckt 4818_7440420039_3.9u 1 2
Rp 1 2 4853
Cp 1 2 1.3p
Rs 1 N3 0.06
L1 N3 2 3.9u
.ends 4818_7440420039_3.9u
*******
.subckt 4818_744042004_4.7u 1 2
Rp 1 2 5535
Cp 1 2 1.24p
Rs 1 N3 0.07
L1 N3 2 4.7u
.ends 4818_744042004_4.7u
*******
.subckt 4818_744042005_5.6u 1 2
Rp 1 2 6390
Cp 1 2 1.42p
Rs 1 N3 0.08
L1 N3 2 5.6u
.ends 4818_744042005_5.6u
*******
.subckt 4818_744042006_6.8u 1 2
Rp 1 2 6793
Cp 1 2 1.51p
Rs 1 N3 0.08
L1 N3 2 6.8u
.ends 4818_744042006_6.8u
*******
.subckt 4818_744042008_8.2u 1 2
Rp 1 2 8512
Cp 1 2 1.54p
Rs 1 N3 0.1
L1 N3 2 8.2u
.ends 4818_744042008_8.2u
*******
.subckt 4818_744042100_10u 1 2
Rp 1 2 10187
Cp 1 2 1.57p
Rs 1 N3 0.12
L1 N3 2 10u
.ends 4818_744042100_10u
*******
.subckt 4818_744042101_100u 1 2
Rp 1 2 36374
Cp 1 2 1.74p
Rs 1 N3 1.17
L1 N3 2 100u
.ends 4818_744042101_100u
*******
.subckt 4818_744042120_12u 1 2
Rp 1 2 10430
Cp 1 2 1.69p
Rs 1 N3 0.15
L1 N3 2 12u
.ends 4818_744042120_12u
*******
.subckt 4818_744042150_15u 1 2
Rp 1 2 13100
Cp 1 2 1.61p
Rs 1 N3 0.19
L1 N3 2 15u
.ends 4818_744042150_15u
*******
.subckt 4818_744042180_18u 1 2
Rp 1 2 14886
Cp 1 2 1.57p
Rs 1 N3 0.27
L1 N3 2 18u
.ends 4818_744042180_18u
*******
.subckt 4818_744042220_22u 1 2
Rp 1 2 16765
Cp 1 2 1.46p
Rs 1 N3 0.28
L1 N3 2 22u
.ends 4818_744042220_22u
*******
.subckt 4818_744042221_220u 1 2
Rp 1 2 54739
Cp 1 2 2.795p
Rs 1 N3 2.88
L1 N3 2 220u
.ends 4818_744042221_220u
*******
.subckt 4818_744042330_33u 1 2
Rp 1 2 18423
Cp 1 2 1.84p
Rs 1 N3 0.382
L1 N3 2 33u
.ends 4818_744042330_33u
*******
.subckt 4818_744042331_330u 1 2
Rp 1 2 85477
Cp 1 2 2.751p
Rs 1 N3 4.1
L1 N3 2 330u
.ends 4818_744042331_330u
*******
.subckt 4818_744042470_47u 1 2
Rp 1 2 20855
Cp 1 2 2.699p
Rs 1 N3 0.54
L1 N3 2 47u
.ends 4818_744042470_47u
*******
.subckt 4818_744042680_68u 1 2
Rp 1 2 27915
Cp 1 2 2.717p
Rs 1 N3 0.715
L1 N3 2 68u
.ends 4818_744042680_68u
*******
.subckt 4828_74404300033_0.33u 1 2
Rp 1 2 385
Cp 1 2 0.489p
Rs 1 N3 0.008
L1 N3 2 0.33u
.ends 4828_74404300033_0.33u
*******
.subckt 4828_74404300047_0.47u 1 2
Rp 1 2 617
Cp 1 2 0.665p
Rs 1 N3 0.01
L1 N3 2 0.47u
.ends 4828_74404300047_0.47u
*******
.subckt 4828_74404300082_0.82u 1 2
Rp 1 2 1023
Cp 1 2 0.795p
Rs 1 N3 0.014
L1 N3 2 0.82u
.ends 4828_74404300082_0.82u
*******
.subckt 4828_7440430012_1.2u 1 2
Rp 1 2 1461
Cp 1 2 0.573p
Rs 1 N3 0.015
L1 N3 2 1.2u
.ends 4828_7440430012_1.2u
*******
.subckt 4828_7440430018_1.8u 1 2
Rp 1 2 1877
Cp 1 2 1.03p
Rs 1 N3 0.02
L1 N3 2 1.8u
.ends 4828_7440430018_1.8u
*******
.subckt 4828_7440430022_2.2u 1 2
Rp 1 2 2395
Cp 1 2 1.33p
Rs 1 N3 0.027
L1 N3 2 2.2u
.ends 4828_7440430022_2.2u
*******
.subckt 4828_7440430027_2.7u 1 2
Rp 1 2 2914
Cp 1 2 1.38p
Rs 1 N3 0.025
L1 N3 2 2.7u
.ends 4828_7440430027_2.7u
*******
.subckt 4828_744043003_3.3u 1 2
Rp 1 2 3425
Cp 1 2 2.16p
Rs 1 N3 0.03
L1 N3 2 3.3u
.ends 4828_744043003_3.3u
*******
.subckt 4828_7440430039_3.9u 1 2
Rp 1 2 2688
Cp 1 2 2.235p
Rs 1 N3 0.05
L1 N3 2 3.9u
.ends 4828_7440430039_3.9u
*******
.subckt 4828_744043004_4.7u 1 2
Rp 1 2 4095
Cp 1 2 1.68p
Rs 1 N3 0.05
L1 N3 2 4.7u
.ends 4828_744043004_4.7u
*******
.subckt 4828_744043005_5.6u 1 2
Rp 1 2 4813
Cp 1 2 0.82p
Rs 1 N3 0.07
L1 N3 2 5.6u
.ends 4828_744043005_5.6u
*******
.subckt 4828_744043006_6.8u 1 2
Rp 1 2 5581
Cp 1 2 1.23p
Rs 1 N3 0.08
L1 N3 2 6.8u
.ends 4828_744043006_6.8u
*******
.subckt 4828_744043008_8.2u 1 2
Rp 1 2 6763
Cp 1 2 1.69p
Rs 1 N3 0.09
L1 N3 2 8.2u
.ends 4828_744043008_8.2u
*******
.subckt 4828_744043100_10u 1 2
Rp 1 2 6973
Cp 1 2 1.944p
Rs 1 N3 0.095
L1 N3 2 10u
.ends 4828_744043100_10u
*******
.subckt 4828_744043101_100u 1 2
Rp 1 2 33813
Cp 1 2 2.94p
Rs 1 N3 0.55
L1 N3 2 100u
.ends 4828_744043101_100u
*******
.subckt 4828_744043102_1000u 1 2
Rp 1 2 180588
Cp 1 2 4.863p
Rs 1 N3 5.4
L1 N3 2 1000u
.ends 4828_744043102_1000u
*******
.subckt 4828_744043120_12u 1 2
Rp 1 2 7529
Cp 1 2 3.36p
Rs 1 N3 0.1
L1 N3 2 12u
.ends 4828_744043120_12u
*******
.subckt 4828_744043150_15u 1 2
Rp 1 2 9705
Cp 1 2 2.65p
Rs 1 N3 0.12
L1 N3 2 15u
.ends 4828_744043150_15u
*******
.subckt 4828_744043151_150u 1 2
Rp 1 2 29583
Cp 1 2 3.55p
Rs 1 N3 0.77
L1 N3 2 150u
.ends 4828_744043151_150u
*******
.subckt 4828_744043152_1500u 1 2
Rp 1 2 103878
Cp 1 2 3.7p
Rs 1 N3 6.8
L1 N3 2 1500u
.ends 4828_744043152_1500u
*******
.subckt 4828_744043180_18u 1 2
Rp 1 2 10720
Cp 1 2 2.38p
Rs 1 N3 0.15
L1 N3 2 18u
.ends 4828_744043180_18u
*******
.subckt 4828_744043220_22u 1 2
Rp 1 2 12152
Cp 1 2 2.44p
Rs 1 N3 0.16
L1 N3 2 22u
.ends 4828_744043220_22u
*******
.subckt 4828_744043221_220u 1 2
Rp 1 2 36973
Cp 1 2 3.55p
Rs 1 N3 1.008
L1 N3 2 220u
.ends 4828_744043221_220u
*******
.subckt 4828_744043270_27u 1 2
Rp 1 2 11258
Cp 1 2 4.339p
Rs 1 N3 0.17
L1 N3 2 27u
.ends 4828_744043270_27u
*******
.subckt 4828_744043330_33u 1 2
Rp 1 2 14941
Cp 1 2 2.81p
Rs 1 N3 0.195
L1 N3 2 33u
.ends 4828_744043330_33u
*******
.subckt 4828_744043331_330u 1 2
Rp 1 2 72822
Cp 1 2 4.292p
Rs 1 N3 1.63
L1 N3 2 330u
.ends 4828_744043331_330u
*******
.subckt 4828_744043390_39u 1 2
Rp 1 2 15149
Cp 1 2 4.228p
Rs 1 N3 0.215
L1 N3 2 39u
.ends 4828_744043390_39u
*******
.subckt 4828_744043470_47u 1 2
Rp 1 2 16524
Cp 1 2 3.39p
Rs 1 N3 0.25
L1 N3 2 47u
.ends 4828_744043470_47u
*******
.subckt 4828_744043471_470u 1 2
Rp 1 2 35458
Cp 1 2 3.6p
Rs 1 N3 2.128
L1 N3 2 470u
.ends 4828_744043471_470u
*******
.subckt 4828_744043561_560u 1 2
Rp 1 2 90660
Cp 1 2 4.619p
Rs 1 N3 2.61
L1 N3 2 560u
.ends 4828_744043561_560u
*******
.subckt 4828_744043680_68u 1 2
Rp 1 2 24607
Cp 1 2 3.12p
Rs 1 N3 0.34
L1 N3 2 68u
.ends 4828_744043680_68u
*******
.subckt 5818_7440520012_1.2u 1 2
Rp 1 2 1478
Cp 1 2 1.26p
Rs 1 N3 0.02
L1 N3 2 1.2u
.ends 5818_7440520012_1.2u
*******
.subckt 5818_7440520018_1.8u 1 2
Rp 1 2 2283
Cp 1 2 1.22p
Rs 1 N3 0.03
L1 N3 2 1.8u
.ends 5818_7440520018_1.8u
*******
.subckt 5818_744052002_2.5u 1 2
Rp 1 2 2612
Cp 1 2 1.66p
Rs 1 N3 0.02
L1 N3 2 2.5u
.ends 5818_744052002_2.5u
*******
.subckt 5818_744052003_3u 1 2
Rp 1 2 3053
Cp 1 2 1.56p
Rs 1 N3 0.04
L1 N3 2 3u
.ends 5818_744052003_3u
*******
.subckt 5818_7440520039_3.9u 1 2
Rp 1 2 4000
Cp 1 2 1.63p
Rs 1 N3 0.05
L1 N3 2 3.9u
.ends 5818_7440520039_3.9u
*******
.subckt 5818_744052005_5u 1 2
Rp 1 2 5060
Cp 1 2 1.7p
Rs 1 N3 0.05
L1 N3 2 5u
.ends 5818_744052005_5u
*******
.subckt 5818_744052006_6.2u 1 2
Rp 1 2 5630
Cp 1 2 1.64p
Rs 1 N3 0.07
L1 N3 2 6.2u
.ends 5818_744052006_6.2u
*******
.subckt 5818_744052007_7.5u 1 2
Rp 1 2 6785
Cp 1 2 1.95p
Rs 1 N3 0.07
L1 N3 2 7.5u
.ends 5818_744052007_7.5u
*******
.subckt 5818_744052009_9u 1 2
Rp 1 2 6970
Cp 1 2 1.72p
Rs 1 N3 0.09
L1 N3 2 9u
.ends 5818_744052009_9u
*******
.subckt 5818_744052100_10u 1 2
Rp 1 2 8291
Cp 1 2 1.68p
Rs 1 N3 0.105
L1 N3 2 10u
.ends 5818_744052100_10u
*******
.subckt 5818_744052101_100u 1 2
Rp 1 2 29220
Cp 1 2 2.735p
Rs 1 N3 0.815
L1 N3 2 100u
.ends 5818_744052101_100u
*******
.subckt 5818_744052120_12u 1 2
Rp 1 2 9612
Cp 1 2 1.57p
Rs 1 N3 0.13
L1 N3 2 12u
.ends 5818_744052120_12u
*******
.subckt 5818_744052150_15u 1 2
Rp 1 2 11201
Cp 1 2 1.29p
Rs 1 N3 0.175
L1 N3 2 15u
.ends 5818_744052150_15u
*******
.subckt 5818_744052180_18u 1 2
Rp 1 2 13516
Cp 1 2 1.64p
Rs 1 N3 0.185
L1 N3 2 18u
.ends 5818_744052180_18u
*******
.subckt 5818_744052220_22u 1 2
Rp 1 2 14029
Cp 1 2 1.6p
Rs 1 N3 0.24
L1 N3 2 22u
.ends 5818_744052220_22u
*******
.subckt 5818_744052221_220u 1 2
Rp 1 2 61323
Cp 1 2 2.195p
Rs 1 N3 2.4
L1 N3 2 220u
.ends 5818_744052221_220u
*******
.subckt 5818_744052270_27u 1 2
Rp 1 2 14180.2
Cp 1 2 1.43p
Rs 1 N3 0.25
L1 N3 2 27u
.ends 5818_744052270_27u
*******
.subckt 5818_744052470_47u 1 2
Rp 1 2 22464
Cp 1 2 1.67p
Rs 1 N3 0.53
L1 N3 2 47u
.ends 5818_744052470_47u
*******
.subckt 5818_744052471_470u 1 2
Rp 1 2 104768
Cp 1 2 2.346p
Rs 1 N3 4.175
L1 N3 2 470u
.ends 5818_744052471_470u
*******
.subckt 5818_744052680_68u 1 2
Rp 1 2 29145
Cp 1 2 1.94p
Rs 1 N3 0.84
L1 N3 2 68u
.ends 5818_744052680_68u
*******
.subckt 5828_744053002_2.6u 1 2
Rp 1 2 2100
Cp 1 2 1.32p
Rs 1 N3 0.02
L1 N3 2 2.6u
.ends 5828_744053002_2.6u
*******
.subckt 5828_744053003_3u 1 2
Rp 1 2 2341
Cp 1 2 2.96p
Rs 1 N3 0.02
L1 N3 2 3u
.ends 5828_744053003_3u
*******
.subckt 5828_744053004_4.2u 1 2
Rp 1 2 2617
Cp 1 2 1.86p
Rs 1 N3 0.03
L1 N3 2 4.2u
.ends 5828_744053004_4.2u
*******
.subckt 5828_7440530047_4.7u 1 2
Rp 1 2 3179
Cp 1 2 2.3p
Rs 1 N3 0.03
L1 N3 2 4.7u
.ends 5828_7440530047_4.7u
*******
.subckt 5828_744053005_5.3u 1 2
Rp 1 2 3981
Cp 1 2 2.24p
Rs 1 N3 0.03
L1 N3 2 5.3u
.ends 5828_744053005_5.3u
*******
.subckt 5828_744053006_6.2u 1 2
Rp 1 2 4071
Cp 1 2 2.2p
Rs 1 N3 0.04
L1 N3 2 6.2u
.ends 5828_744053006_6.2u
*******
.subckt 5828_744053008_8.2u 1 2
Rp 1 2 6785
Cp 1 2 1.95p
Rs 1 N3 0.05
L1 N3 2 8.2u
.ends 5828_744053008_8.2u
*******
.subckt 5828_744053100_10u 1 2
Rp 1 2 6970
Cp 1 2 1.72p
Rs 1 N3 0.06
L1 N3 2 10u
.ends 5828_744053100_10u
*******
.subckt 5828_744053101_100u 1 2
Rp 1 2 24206
Cp 1 2 3.11p
Rs 1 N3 0.4
L1 N3 2 100u
.ends 5828_744053101_100u
*******
.subckt 5828_744053120_12u 1 2
Rp 1 2 6728
Cp 1 2 3.63p
Rs 1 N3 0.07
L1 N3 2 12u
.ends 5828_744053120_12u
*******
.subckt 5828_744053150_15u 1 2
Rp 1 2 6970
Cp 1 2 2.9p
Rs 1 N3 0.08
L1 N3 2 15u
.ends 5828_744053150_15u
*******
.subckt 5828_744053180_18u 1 2
Rp 1 2 9311
Cp 1 2 3.6p
Rs 1 N3 0.09
L1 N3 2 18u
.ends 5828_744053180_18u
*******
.subckt 5828_744053220_22u 1 2
Rp 1 2 9672
Cp 1 2 2.76p
Rs 1 N3 0.1
L1 N3 2 22u
.ends 5828_744053220_22u
*******
.subckt 5828_744053221_220u 1 2
Rp 1 2 61323
Cp 1 2 2.19p
Rs 1 N3 1.17
L1 N3 2 220u
.ends 5828_744053221_220u
*******
.subckt 5828_744053270_27u 1 2
Rp 1 2 13015
Cp 1 2 2.85p
Rs 1 N3 0.135
L1 N3 2 27u
.ends 5828_744053270_27u
*******
.subckt 5828_744053330_33u 1 2
Rp 1 2 13481
Cp 1 2 2.89p
Rs 1 N3 0.18
L1 N3 2 33u
.ends 5828_744053330_33u
*******
.subckt 5828_744053470_47u 1 2
Rp 1 2 18925
Cp 1 2 3.07p
Rs 1 N3 0.22
L1 N3 2 47u
.ends 5828_744053470_47u
*******
.subckt 5828_744053680_68u 1 2
Rp 1 2 24200
Cp 1 2 2.79p
Rs 1 N3 0.3
L1 N3 2 68u
.ends 5828_744053680_68u
*******
.subckt 6823_744062001_1u 1 2
Rp 1 2 883
Cp 1 2 1.28p
Rs 1 N3 0.01
L1 N3 2 1u
.ends 6823_744062001_1u
*******
.subckt 6823_7440620015_1.5u 1 2
Rp 1 2 1383
Cp 1 2 1.63p
Rs 1 N3 0.01
L1 N3 2 1.5u
.ends 6823_7440620015_1.5u
*******
.subckt 6823_744062002_2.2u 1 2
Rp 1 2 2019
Cp 1 2 2.03p
Rs 1 N3 0.01
L1 N3 2 2.2u
.ends 6823_744062002_2.2u
*******
.subckt 6823_744062003_3.3u 1 2
Rp 1 2 2700
Cp 1 2 2.28p
Rs 1 N3 0.02
L1 N3 2 3.3u
.ends 6823_744062003_3.3u
*******
.subckt 6823_744062005_5u 1 2
Rp 1 2 3361
Cp 1 2 2.03p
Rs 1 N3 0.04
L1 N3 2 5u
.ends 6823_744062005_5u
*******
.subckt 6823_744062006_6.2u 1 2
Rp 1 2 4645
Cp 1 2 2.44p
Rs 1 N3 0.04
L1 N3 2 6.2u
.ends 6823_744062006_6.2u
*******
.subckt 6823_744062007_7.5u 1 2
Rp 1 2 5466
Cp 1 2 2.14p
Rs 1 N3 0.05
L1 N3 2 7.5u
.ends 6823_744062007_7.5u
*******
.subckt 6823_744062100_10u 1 2
Rp 1 2 6728
Cp 1 2 2.04p
Rs 1 N3 0.053
L1 N3 2 10u
.ends 6823_744062100_10u
*******
.subckt 6823_744062101_100u 1 2
Rp 1 2 32358
Cp 1 2 2.48p
Rs 1 N3 0.44
L1 N3 2 100u
.ends 6823_744062101_100u
*******
.subckt 6823_744062102_1000u 1 2
Rp 1 2 109964
Cp 1 2 3.11p
Rs 1 N3 3.82
L1 N3 2 1000u
.ends 6823_744062102_1000u
*******
.subckt 6823_744062120_12u 1 2
Rp 1 2 5990
Cp 1 2 2.41p
Rs 1 N3 0.07
L1 N3 2 12u
.ends 6823_744062120_12u
*******
.subckt 6823_744062150_15u 1 2
Rp 1 2 9100
Cp 1 2 2.48p
Rs 1 N3 0.08
L1 N3 2 15u
.ends 6823_744062150_15u
*******
.subckt 6823_744062151_150u 1 2
Rp 1 2 53810
Cp 1 2 2.37p
Rs 1 N3 0.605
L1 N3 2 150u
.ends 6823_744062151_150u
*******
.subckt 6823_744062152_1500u 1 2
Rp 1 2 187958
Cp 1 2 2.66p
Rs 1 N3 7
L1 N3 2 1500u
.ends 6823_744062152_1500u
*******
.subckt 6823_744062180_18u 1 2
Rp 1 2 8675
Cp 1 2 2.28p
Rs 1 N3 0.09
L1 N3 2 18u
.ends 6823_744062180_18u
*******
.subckt 6823_744062220_22u 1 2
Rp 1 2 10662
Cp 1 2 2.42p
Rs 1 N3 0.1
L1 N3 2 22u
.ends 6823_744062220_22u
*******
.subckt 6823_744062221_220u 1 2
Rp 1 2 61452.5
Cp 1 2 1.971p
Rs 1 N3 1.01
L1 N3 2 220u
.ends 6823_744062221_220u
*******
.subckt 6823_744062330_33u 1 2
Rp 1 2 17164
Cp 1 2 2.16p
Rs 1 N3 0.15
L1 N3 2 33u
.ends 6823_744062330_33u
*******
.subckt 6823_744062470_47u 1 2
Rp 1 2 19143
Cp 1 2 2.96p
Rs 1 N3 0.26
L1 N3 2 47u
.ends 6823_744062470_47u
*******
.subckt 6823_744062680_68u 1 2
Rp 1 2 23150
Cp 1 2 2.27p
Rs 1 N3 0.3
L1 N3 2 68u
.ends 6823_744062680_68u
*******
.subckt 8012_74406800024_0.24u 1 2
Rp 1 2 338
Cp 1 2 0.187p
Rs 1 N3 0.015
L1 N3 2 0.24u
.ends 8012_74406800024_0.24u
*******
.subckt 8012_74406800056_0.56u 1 2
Rp 1 2 813
Cp 1 2 0.541p
Rs 1 N3 0.022
L1 N3 2 0.56u
.ends 8012_74406800056_0.56u
*******
.subckt 8012_7440680010_1u 1 2
Rp 1 2 1500
Cp 1 2 0.924p
Rs 1 N3 0.032
L1 N3 2 1u
.ends 8012_7440680010_1u
*******
.subckt 8012_7440680017_1.7u 1 2
Rp 1 2 2132
Cp 1 2 1.36p
Rs 1 N3 0.041
L1 N3 2 1.7u
.ends 8012_7440680017_1.7u
*******
.subckt 8012_7440680027_2.7u 1 2
Rp 1 2 2856
Cp 1 2 1.57p
Rs 1 N3 0.052
L1 N3 2 2.7u
.ends 8012_7440680027_2.7u
*******
.subckt 8012_7440680033_3.3u 1 2
Rp 1 2 3804
Cp 1 2 1.73p
Rs 1 N3 0.061
L1 N3 2 3.3u
.ends 8012_7440680033_3.3u
*******
.subckt 8012_7440680047_4.7u 1 2
Rp 1 2 4377
Cp 1 2 1.95p
Rs 1 N3 0.072
L1 N3 2 4.7u
.ends 8012_7440680047_4.7u
*******
.subckt 8012_7440680056_5.6u 1 2
Rp 1 2 6305
Cp 1 2 1.43p
Rs 1 N3 0.11
L1 N3 2 5.6u
.ends 8012_7440680056_5.6u
*******
.subckt 8012_7440680068_6.8u 1 2
Rp 1 2 6807
Cp 1 2 1.71p
Rs 1 N3 0.127
L1 N3 2 6.8u
.ends 8012_7440680068_6.8u
*******
.subckt 8012_7440680082_8.2u 1 2
Rp 1 2 7101
Cp 1 2 1.52p
Rs 1 N3 0.142
L1 N3 2 8.2u
.ends 8012_7440680082_8.2u
*******
.subckt 8012_7440680100_10u 1 2
Rp 1 2 8000
Cp 1 2 2.32p
Rs 1 N3 0.177
L1 N3 2 10u
.ends 8012_7440680100_10u
*******
.subckt 8012_7440680120_12u 1 2
Rp 1 2 9131
Cp 1 2 2.31p
Rs 1 N3 0.195
L1 N3 2 12u
.ends 8012_7440680120_12u
*******
.subckt 8012_7440680150_15u 1 2
Rp 1 2 8188
Cp 1 2 3.18p
Rs 1 N3 0.213
L1 N3 2 15u
.ends 8012_7440680150_15u
*******
.subckt 8012_7440680180_18u 1 2
Rp 1 2 10907
Cp 1 2 3.02p
Rs 1 N3 0.302
L1 N3 2 18u
.ends 8012_7440680180_18u
*******
.subckt 8012_7440680220_22u 1 2
Rp 1 2 11969
Cp 1 2 3.49p
Rs 1 N3 0.35
L1 N3 2 22u
.ends 8012_7440680220_22u
*******
.subckt 8015_74406900022_0.22u 1 2
Rp 1 2 330
Cp 1 2 0.177p
Rs 1 N3 0.009
L1 N3 2 0.22u
.ends 8015_74406900022_0.22u
*******
.subckt 8015_74406900052_0.52u 1 2
Rp 1 2 780
Cp 1 2 0.5p
Rs 1 N3 0.015
L1 N3 2 0.52u
.ends 8015_74406900052_0.52u
*******
.subckt 8015_7440690010_1u 1 2
Rp 1 2 1445
Cp 1 2 0.65p
Rs 1 N3 0.021
L1 N3 2 1u
.ends 8015_7440690010_1u
*******
.subckt 8015_7440690016_1.6u 1 2
Rp 1 2 2240
Cp 1 2 0.82p
Rs 1 N3 0.029
L1 N3 2 1.6u
.ends 8015_7440690016_1.6u
*******
.subckt 8015_7440690022_2.2u 1 2
Rp 1 2 3222
Cp 1 2 1.07p
Rs 1 N3 0.035
L1 N3 2 2.2u
.ends 8015_7440690022_2.2u
*******
.subckt 8015_7440690033_3.3u 1 2
Rp 1 2 3803
Cp 1 2 1.34p
Rs 1 N3 0.042
L1 N3 2 3.3u
.ends 8015_7440690033_3.3u
*******
.subckt 8015_7440690047_4.7u 1 2
Rp 1 2 4853
Cp 1 2 1.33p
Rs 1 N3 0.056
L1 N3 2 4.7u
.ends 8015_7440690047_4.7u
*******
.subckt 8015_7440690068_6.8u 1 2
Rp 1 2 7277
Cp 1 2 1.71p
Rs 1 N3 0.088
L1 N3 2 6.8u
.ends 8015_7440690068_6.8u
*******
.subckt 8015_7440690082_8.2u 1 2
Rp 1 2 8123
Cp 1 2 2.04p
Rs 1 N3 0.099
L1 N3 2 8.2u
.ends 8015_7440690082_8.2u
*******
.subckt 8015_7440690100_10u 1 2
Rp 1 2 7700
Cp 1 2 2.43p
Rs 1 N3 0.112
L1 N3 2 10u
.ends 8015_7440690100_10u
*******
.subckt 8015_7440690120_12u 1 2
Rp 1 2 9407
Cp 1 2 2.13p
Rs 1 N3 0.148
L1 N3 2 12u
.ends 8015_7440690120_12u
*******
.subckt 8015_7440690150_15u 1 2
Rp 1 2 11103
Cp 1 2 2.75p
Rs 1 N3 0.179
L1 N3 2 15u
.ends 8015_7440690150_15u
*******
.subckt 8015_7440690180_18u 1 2
Rp 1 2 13318
Cp 1 2 3.03p
Rs 1 N3 0.225
L1 N3 2 18u
.ends 8015_7440690180_18u
*******
.subckt 8015_7440690220_22u 1 2
Rp 1 2 14590
Cp 1 2 2.68p
Rs 1 N3 0.272
L1 N3 2 22u
.ends 8015_7440690220_22u
*******
.subckt 8020_74407000018_0.18u 1 2
Rp 1 2 290
Cp 1 2 0.633p
Rs 1 N3 0.00351
L1 N3 2 0.18u
.ends 8020_74407000018_0.18u
*******
.subckt 8020_74407000047_0.47u 1 2
Rp 1 2 612
Cp 1 2 1p
Rs 1 N3 0.0058
L1 N3 2 0.47u
.ends 8020_74407000047_0.47u
*******
.subckt 8020_74407000082_0.82u 1 2
Rp 1 2 1006
Cp 1 2 1.455p
Rs 1 N3 0.0085
L1 N3 2 0.82u
.ends 8020_74407000082_0.82u
*******
.subckt 8020_7440700012_1.2u 1 2
Rp 1 2 1680
Cp 1 2 1.56p
Rs 1 N3 0.0125
L1 N3 2 1.2u
.ends 8020_7440700012_1.2u
*******
.subckt 8020_7440700022_2.2u 1 2
Rp 1 2 2000
Cp 1 2 1.88p
Rs 1 N3 0.017
L1 N3 2 2.2u
.ends 8020_7440700022_2.2u
*******
.subckt 8020_7440700033_3.3u 1 2
Rp 1 2 2900
Cp 1 2 2.13p
Rs 1 N3 0.03
L1 N3 2 3.3u
.ends 8020_7440700033_3.3u
*******
.subckt 8020_7440700047_4.7u 1 2
Rp 1 2 3470
Cp 1 2 2p
Rs 1 N3 0.037
L1 N3 2 4.7u
.ends 8020_7440700047_4.7u
*******
.subckt 8020_7440700056_5.6u 1 2
Rp 1 2 4174
Cp 1 2 2.05p
Rs 1 N3 0.047
L1 N3 2 5.6u
.ends 8020_7440700056_5.6u
*******
.subckt 8020_7440700068_6.8u 1 2
Rp 1 2 4000
Cp 1 2 2.1p
Rs 1 N3 0.056
L1 N3 2 6.8u
.ends 8020_7440700068_6.8u
*******
.subckt 8020_7440700082_8.2u 1 2
Rp 1 2 5120
Cp 1 2 2.1p
Rs 1 N3 0.0705
L1 N3 2 8.2u
.ends 8020_7440700082_8.2u
*******
.subckt 8020_7440700100_10u 1 2
Rp 1 2 5500
Cp 1 2 2.17p
Rs 1 N3 0.078
L1 N3 2 10u
.ends 8020_7440700100_10u
*******
.subckt 8020_7440700150_15u 1 2
Rp 1 2 6900
Cp 1 2 2.26p
Rs 1 N3 0.117
L1 N3 2 15u
.ends 8020_7440700150_15u
*******
.subckt 8020_7440700180_18u 1 2
Rp 1 2 7520
Cp 1 2 2.4p
Rs 1 N3 0.135
L1 N3 2 18u
.ends 8020_7440700180_18u
*******
.subckt 8020_7440700220_22u 1 2
Rp 1 2 9000
Cp 1 2 2.4p
Rs 1 N3 0.166
L1 N3 2 22u
.ends 8020_7440700220_22u
*******
.subckt 8043_7440710082_0.82u 1 2
Rp 1 2 1174
Cp 1 2 2.3321p
Rs 1 N3 0.007
L1 N3 2 0.82u
.ends 8043_7440710082_0.82u
*******
.subckt 8043_744071022_2.2u 1 2
Rp 1 2 2730
Cp 1 2 3.92p
Rs 1 N3 0.01
L1 N3 2 2.2u
.ends 8043_744071022_2.2u
*******
.subckt 8043_744071039_3.9u 1 2
Rp 1 2 4061
Cp 1 2 4.58p
Rs 1 N3 0.013
L1 N3 2 3.9u
.ends 8043_744071039_3.9u
*******
.subckt 8043_744071047_4.7u 1 2
Rp 1 2 4986
Cp 1 2 4.34p
Rs 1 N3 0.017
L1 N3 2 4.7u
.ends 8043_744071047_4.7u
*******
.subckt 8043_744071056_5.6u 1 2
Rp 1 2 5843
Cp 1 2 5.05p
Rs 1 N3 0.02
L1 N3 2 5.6u
.ends 8043_744071056_5.6u
*******
.subckt 8043_744071100_10u 1 2
Rp 1 2 7595
Cp 1 2 5.32p
Rs 1 N3 0.028
L1 N3 2 10u
.ends 8043_744071100_10u
*******
.subckt 8043_744071101_100u 1 2
Rp 1 2 67323
Cp 1 2 6.8p
Rs 1 N3 0.27
L1 N3 2 100u
.ends 8043_744071101_100u
*******
.subckt 8043_744071102_1m 1 2
Rp 1 2 349863
Cp 1 2 6.11p
Rs 1 N3 2.985
L1 N3 2 1000u
.ends 8043_744071102_1m
*******
.subckt 8043_744071150_15u 1 2
Rp 1 2 12488
Cp 1 2 5.02p
Rs 1 N3 0.046
L1 N3 2 15u
.ends 8043_744071150_15u
*******
.subckt 8043_744071220_22u 1 2
Rp 1 2 14321
Cp 1 2 5.09p
Rs 1 N3 0.065
L1 N3 2 22u
.ends 8043_744071220_22u
*******
.subckt 8043_744071221_220u 1 2
Rp 1 2 94497
Cp 1 2 5.885p
Rs 1 N3 0.51
L1 N3 2 220u
.ends 8043_744071221_220u
*******
.subckt 8043_744071330_33u 1 2
Rp 1 2 18901
Cp 1 2 5.56p
Rs 1 N3 0.095
L1 N3 2 33u
.ends 8043_744071330_33u
*******
.subckt 8043_744071470_47u 1 2
Rp 1 2 28491
Cp 1 2 5.82p
Rs 1 N3 0.12
L1 N3 2 47u
.ends 8043_744071470_47u
*******
.subckt 8043_744071680_68u 1 2
Rp 1 2 35800
Cp 1 2 6.81p
Rs 1 N3 0.185
L1 N3 2 68u
.ends 8043_744071680_68u
*******
