**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT High Current Inductor
* Matchcode:             WE-CHSA
* Library Type:          LTspice
* Version:               rev21a
* Created/modified by:   Ella
* Date and Time:         2022/10/27
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
.subckt 1011_7843330033_0.33u 1 2
Rp 1 2 173.347
Cp 1 2 1.5p
Rs 1 N3 0.0014
L1 N3 2 0.350437u
.ends 1011_7843330033_0.33u
*******
.subckt 1011_7843330056_0.56u 1 2
Rp 1 2 327.941
Cp 1 2 4.14p
Rs 1 N3 0.0017
L1 N3 2 0.611835u
.ends 1011_7843330056_0.56u
*******
.subckt 1011_7843330100_1u 1 2
Rp 1 2 538.519
Cp 1 2 3.416p
Rs 1 N3 0.0024
L1 N3 2 0.915553u
.ends 1011_7843330100_1u
*******
.subckt 1011_7843330180_1.8u 1 2
Rp 1 2 1113
Cp 1 2 3.38p
Rs 1 N3 0.0039
L1 N3 2 1.783u
.ends 1011_7843330180_1.8u
*******
.subckt 1011_7843330330_3.3u 1 2
Rp 1 2 1872
Cp 1 2 2.769p
Rs 1 N3 0.0054
L1 N3 2 2.958u
.ends 1011_7843330330_3.3u
*******
.subckt 1011_7843330390_3.9u 1 2
Rp 1 2 2228
Cp 1 2 2.4846733735p
Rs 1 N3 0.00725
L1 N3 2 3.406u
.ends 1011_7843330390_3.9u
*******
.subckt 1011_7843330560_5.6u 1 2
Rp 1 2 3691
Cp 1 2 3.017p
Rs 1 N3 0.01085
L1 N3 2 5.297u
.ends 1011_7843330560_5.6u
*******
.subckt 1011_7843330820_8.2u 1 2
Rp 1 2 4914
Cp 1 2 3.221p
Rs 1 N3 0.0159
L1 N3 2 6.921u
.ends 1011_7843330820_8.2u
*******
.subckt 1011_7843331000_10u 1 2
Rp 1 2 5588
Cp 1 2 3.239p
Rs 1 N3 0.0215
L1 N3 2 8.652u
.ends 1011_7843331000_10u
*******
.subckt 1011_7843331200_12u 1 2
Rp 1 2 9806.78338388
Cp 1 2 2.42581600528p
Rs 1 N3 0.0277
L1 N3 2 12.6279218099u
.ends 1011_7843331200_12u
*******
.subckt 1011_7843331800_18u 1 2
Rp 1 2 12350
Cp 1 2 2.922p
Rs 1 N3 0.03425
L1 N3 2 15.888u
.ends 1011_7843331800_18u
*******
.subckt 1011_7843332000_20u 1 2
Rp 1 2 13884
Cp 1 2 2.917p
Rs 1 N3 0.0508
L1 N3 2 20.163u
.ends 1011_7843332000_20u
*******
.subckt 1212_7843320039_0.39u 1 2
Rp 1 2 161.175
Cp 1 2 7.28p
Rs 1 N3 0.00135
L1 N3 2 0.348075u
.ends 1212_7843320039_0.39u
*******
.subckt 1212_7843320068_0.68u 1 2
Rp 1 2 289.234
Cp 1 2 5.6p
Rs 1 N3 0.0017
L1 N3 2 0.579173u
.ends 1212_7843320068_0.68u
*******
.subckt 1212_7843320100_1u 1 2
Rp 1 2 482.699
Cp 1 2 3.85p
Rs 1 N3 0.002
L1 N3 2 1.001u
.ends 1212_7843320100_1u
*******
.subckt 1212_7843320150_1.5u 1 2
Rp 1 2 853.40702436469
Cp 1 2 2.91228430955172p
Rs 1 N3 0.0027
L1 N3 2 1.55489890604933u
.ends 1212_7843320150_1.5u
*******
.subckt 1212_7843320270_2.7u 1 2
Rp 1 2 1380
Cp 1 2 4.1p
Rs 1 N3 0.0039
L1 N3 2 2.478u
.ends 1212_7843320270_2.7u
*******
.subckt 1212_7843320330_3.3u 1 2
Rp 1 2 1256
Cp 1 2 3.7p
Rs 1 N3 0.0053
L1 N3 2 3.396u
.ends 1212_7843320330_3.3u
*******
.subckt 1212_7843320470_4.7u 1 2
Rp 1 2 2719
Cp 1 2 3.639p
Rs 1 N3 0.00685
L1 N3 2 4.928u
.ends 1212_7843320470_4.7u
*******
.subckt 1212_7843320680_6.8u 1 2
Rp 1 2 3982
Cp 1 2 2.75p
Rs 1 N3 0.0099
L1 N3 2 6.703u
.ends 1212_7843320680_6.8u
*******
.subckt 1212_7843320820_8.2u 1 2
Rp 1 2 4871
Cp 1 2 3.553p
Rs 1 N3 0.01245
L1 N3 2 7.887u
.ends 1212_7843320820_8.2u
*******
.subckt 1212_7843321000_10u 1 2
Rp 1 2 5243
Cp 1 2 3.22p
Rs 1 N3 0.01695
L1 N3 2 8.7u
.ends 1212_7843321000_10u
*******
.subckt 1212_7843321200_12u 1 2
Rp 1 2 7227.97
Cp 1 2 2.83341268310714p
Rs 1 N3 0.0179
L1 N3 2 10.7689388817107u
.ends 1212_7843321200_12u
*******
.subckt 1212_7843321800_18u 1 2
Rp 1 2 11674.8658463
Cp 1 2 3.30968658028p
Rs 1 N3 0.032
L1 N3 2 17.4350688226u
.ends 1212_7843321800_18u
*******
.subckt 1212_7843322000_20u 1 2
Rp 1 2 14544
Cp 1 2 3.664p
Rs 1 N3 0.0359
L1 N3 2 20.227u
.ends 1212_7843322000_20u
*******
.subckt 8090_7843340033_0.33u 1 2
Rp 1 2 289.506
Cp 1 2 2.1p
Rs 1 N3 0.00175
L1 N3 2 0.312059u
.ends 8090_7843340033_0.33u
*******
.subckt 8090_7843340047_0.47u 1 2
Rp 1 2 468.308
Cp 1 2 2.62p
Rs 1 N3 0.0023
L1 N3 2 0.452357u
.ends 8090_7843340047_0.47u
*******
.subckt 8090_7843340068_0.68u 1 2
Rp 1 2 682.666
Cp 1 2 1.94p
Rs 1 N3 0.00345
L1 N3 2 0.746687u
.ends 8090_7843340068_0.68u
*******
.subckt 8090_7843340100_1u 1 2
Rp 1 2 985.376
Cp 1 2 2.45p
Rs 1 N3 0.0049
L1 N3 2 1.028u
.ends 8090_7843340100_1u
*******
.subckt 8090_7843340220_2.2u 1 2
Rp 1 2 2186
Cp 1 2 2.501p
Rs 1 N3 0.01
L1 N3 2 2.24u
.ends 8090_7843340220_2.2u
*******
.subckt 8090_7843340330_3.3u 1 2
Rp 1 2 3271
Cp 1 2 1.7p
Rs 1 N3 0.01535
L1 N3 2 3.287u
.ends 8090_7843340330_3.3u
*******
.subckt 8090_7843340470_4.7u 1 2
Rp 1 2 5206
Cp 1 2 1.994p
Rs 1 N3 0.0241
L1 N3 2 5.057u
.ends 8090_7843340470_4.7u
*******
.subckt 1011_78433390150_1.5u 1 2
Rp 1 2 1602
Cp 1 2 2.823p
Rs 1 N3 0.0039
L1 N3 2 1.388u
.ends 1011_78433390150_1.5u
*******
.subckt 1011_78433390240_2.4u 1 2
Rp 1 2 2607
Cp 1 2 3.048p
Rs 1 N3 0.0054
L1 N3 2 2.278u
.ends 1011_78433390240_2.4u
*******
.subckt 1011_78433390300_3u 1 2
Rp 1 2 3270
Cp 1 2 2.916p
Rs 1 N3 0.00725
L1 N3 2 2.834u
.ends 1011_78433390300_3u
*******
.subckt 1011_78433390430_4.3u 1 2
Rp 1 2 4417
Cp 1 2 3.108p
Rs 1 N3 0.01085
L1 N3 2 4.233u
.ends 1011_78433390430_4.3u
*******
.subckt 1011_78433390620_6.2u 1 2
Rp 1 2 6737
Cp 1 2 2.606p
Rs 1 N3 0.0159
L1 N3 2 5.995u
.ends 1011_78433390620_6.2u
*******
.subckt 1011_78433390820_8.2u 1 2
Rp 1 2 8222
Cp 1 2 3.205p
Rs 1 N3 0.0215
L1 N3 2 7.712u
.ends 1011_78433390820_8.2u
*******
.subckt 1011_78433391000_10u 1 2
Rp 1 2 10415
Cp 1 2 2.911p
Rs 1 N3 0.0277
L1 N3 2 9.504u
.ends 1011_78433391000_10u
*******
.subckt 1011_78433391500_15u 1 2
Rp 1 2 16030
Cp 1 2 3.179p
Rs 1 N3 0.0508
L1 N3 2 15.425u
.ends 1011_78433391500_15u
*******
.subckt 1212_78433290200_2u 1 2
Rp 1 2 1836
Cp 1 2 3.178p
Rs 1 N3 0.0039
L1 N3 2 1.942u
.ends 1212_78433290200_2u
*******
.subckt 1212_78433290240_2.4u 1 2
Rp 1 2 2324
Cp 1 2 2.915p
Rs 1 N3 0.0053
L1 N3 2 2.382u
.ends 1212_78433290240_2.4u
*******
.subckt 1212_78433290360_3.6u 1 2
Rp 1 2 3432
Cp 1 2 3.034p
Rs 1 N3 0.00685
L1 N3 2 3.529u
.ends 1212_78433290360_3.6u
*******
.subckt 1212_78433290510_5.1u 1 2
Rp 1 2 4856
Cp 1 2 2.876p
Rs 1 N3 0.0099
L1 N3 2 5.432u
.ends 1212_78433290510_5.1u
*******
.subckt 1212_78433290620_6.2u 1 2
Rp 1 2 5621
Cp 1 2 3.089p
Rs 1 N3 0.01245
L1 N3 2 6.103u
.ends 1212_78433290620_6.2u
*******
.subckt 1212_78433290750_7.5u 1 2
Rp 1 2 6972
Cp 1 2 2.975p
Rs 1 N3 0.01695
L1 N3 2 7.261u
.ends 1212_78433290750_7.5u
*******
.subckt 1212_78433290820_8.2u 1 2
Rp 1 2 7621
Cp 1 2 3.027p
Rs 1 N3 0.0179
L1 N3 2 8.163u
.ends 1212_78433290820_8.2u
*******
.subckt 1212_78433291500_15u 1 2
Rp 1 2 15563
Cp 1 2 2.89p
Rs 1 N3 0.0359
L1 N3 2 16.066u
.ends 1212_78433291500_15u
*******
.subckt 8090_78433490036_0.36u 1 2
Rp 1 2 751.778
Cp 1 2 1.494p
Rs 1 N3 0.0023
L1 N3 2 0.355435u
.ends 8090_78433490036_0.36u
*******
.subckt 8090_78433490056_0.56u 1 2
Rp 1 2 1078
Cp 1 2 1.449p
Rs 1 N3 0.00345
L1 N3 2 0.514054u
.ends 8090_78433490056_0.56u
*******
.subckt 8090_78433490075_0.75u 1 2
Rp 1 2 1457
Cp 1 2 1.476p
Rs 1 N3 0.0049
L1 N3 2 0.725695u
.ends 8090_78433490075_0.75u
*******
.subckt 8090_78433490160_1.6u 1 2
Rp 1 2 3108
Cp 1 2 1.848p
Rs 1 N3 0.01
L1 N3 2 1.586u
.ends 8090_78433490160_1.6u
*******
.subckt 8090_78433490240_2.4u 1 2
Rp 1 2 4484
Cp 1 2 1.701p
Rs 1 N3 0.01535
L1 N3 2 2.325u
.ends 8090_78433490240_2.4u
*******
.subckt 8090_78433490390_3.9u 1 2
Rp 1 2 6650
Cp 1 2 1.603p
Rs 1 N3 0.0241
L1 N3 2 3.726u
.ends 8090_78433490390_3.9u
*******
