**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Mono-color TOP LED Waterclear
* Matchcode:              WL-SMTW
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-23
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 2214_150224AS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=10.000E-21
+ N=1.7534
+ RS=1.0001E-6
+ IKF=1.8327E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=1.5
+ IBV=5.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224BS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=39.446E-18
+ N=3.0271
+ RS=.99109
+ IKF=182.17E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=1.5
+ IBV=5.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224GS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=47.668E-3
+ N=4.2719
+ RS=3.3656
+ IKF=29.082E-15
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=1.5
+ IBV=5.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224SS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=279.66E-12
+ N=4.3941
+ RS=1.1366
+ IKF=519.47
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=1.5
+ IBV=5.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224YS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=192.98E-12
+ N=4.2946
+ RS=1.0810
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=1.5
+ IBV=5.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224BS73100A  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=16.888E-15
+ N=3.8735
+ RS=1.5380
+ IKF=217.16E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224GS73100A 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=42.238E-12
+ N=4.9113
+ RS=2.6655
+ IKF=307.33E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224RS73100A 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=1.3208E-15
+ N=2.2823
+ RS=.83386
+ IKF=200.04E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224VS73100A 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=635.69E-18
+ N=2.2278
+ RS=.79472
+ IKF=195.42E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2214_150224YS73100A 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=635.69E-18
+ N=2.2278
+ RS=.79472
+ IKF=195.42E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_150283BS73103  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=27.398E-12
+ N=4.5312
+ RS=.24906
+ IKF=1.7137E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_150283GS73103  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=7.5809E-12
+ N=4.0552
+ RS=.21401
+ IKF=1.5730E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_150283RS73103  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=381.17E-12
+ N=4.2460
+ RS=1.0000E-6
+ IKF=.43019
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_150283YS73103 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=588.88E-18
+ N=2.2102
+ RS=88.143E-3
+ IKF=1.0248E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_150283DS73103 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=27.398E-12
+ N=4.5312
+ RS=.24906
+ IKF=1.7137E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_150283FS73103 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=588.88E-18
+ N=2.2102
+ RS=88.143E-3
+ IKF=1.0248E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 2835_150283HS73103 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=588.88E-18
+ N=2.2102
+ RS=88.143E-3
+ IKF=1.0248E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3020_150302BS73100 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=695.94E-6
+ N=5
+ RS=2.4677
+ IKF=16.109E-12
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3020_150302GS73100 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=82.822E-12
+ N=5
+ RS=1.8037
+ IKF=257.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3020_150302RS73100 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=557.55E-18
+ N=2.1602
+ RS=.37378
+ IKF=236.66E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3020_150302VS73100 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=557.55E-18
+ N=2.1602
+ RS=.37378
+ IKF=236.66E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3020_150302YS73100 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=824.78E-18
+ N=2.2038
+ RS=.38595
+ IKF=240.07E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141AS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=557.55E-18
+ N=2.1602
+ RS=.37378
+ IKF=236.66E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141BS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=695.94E-6
+ N=5
+ RS=2.4677
+ IKF=16.109E-12
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141GS73100 1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=2.0835E-6
+ N=4.7862
+ RS=2.1709
+ IKF=3.7697E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141RS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=557.55E-18
+ N=2.1602
+ RS=.37378
+ IKF=236.66E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141VS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=557.55E-18
+ N=2.1602
+ RS=.37378
+ IKF=236.66E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
*****
.subckt 3528_150141YS73100  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=557.55E-18
+ N=2.1602
+ RS=.37378
+ IKF=236.66E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141AS73113 1  2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=26.367E-15
+ N=2.6750
+ RS=.5534
+ IKF=266.68E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141BS73113 1  2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=86.213E-12
+ N=5
+ RS=2.5356
+ IKF=135.10E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141GS73113 1  2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=79.244E-12
+ N=4.9872
+ RS=1.2654
+ IKF=448.72E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141RS73113 1  2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=28.480E-15
+ N=2.6859
+ RS=.52064
+ IKF=276.58E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141YS73113 1  2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=28.480E-15
+ N=2.6859
+ RS=.52064
+ IKF=276.58E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3528_150141BS73130 1 2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=48.651E-12
+ N=4.7513
+ RS=1.1837
+ IKF=431.41E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141BS73140 1 2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=48.651E-12
+ N=4.7513
+ RS=1.1837
+ IKF=431.41E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
***********
.subckt 3528_150141GS73130 1 2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=59.184E-12
+ N=4.8435
+ RS=1.2147
+ IKF=438.32E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141GS73140 1 2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=59.184E-12
+ N=4.8435
+ RS=1.2147
+ IKF=438.32E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
***********
.subckt 3528_150141RS73130 1 2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=201.79E-15
+ N=3.0464
+ RS=.62959
+ IKF=303.48E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141RS73140 1 2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=201.79E-15
+ N=3.0464
+ RS=.62959
+ IKF=303.48E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141YS73130 1 2
D1 1  2 SMTW
.MODEL SMTW D
+ IS=51.276E-15
+ N=2.7856
+ RS=.54975
+ IKF=284.26E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141YS73140 1 2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=51.276E-15
+ N=2.7856
+ RS=.54975
+ IKF=284.26E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
***********
.subckt 5050_150505BS73300  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=76.911E-9
+ N=4.0185
+ RS=1.6401
+ IKF=14.505E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 5050_150505GS73300  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=62.468E-12
+ N=4.8695
+ RS=1.2283
+ IKF=438.14E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 5050_150505RS73300  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=23.817E-18
+ N=1.8613
+ RS=.29697
+ IKF=212.34E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 5050_150505YS73300  1  2
D1 1 2 SMTW
.MODEL SMTW D
+ IS=23.817E-18
+ N=1.8613
+ RS=.29697
+ IKF=212.34E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******





