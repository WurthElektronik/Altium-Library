**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  SMT Power Inductor
* Matchcode:              WE-XHMI
* Library Type:           LTspice
* Version:                rev25b
* Created/modified by:    Ella
* Date and Time:          5/8/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1010P_7443936050022_0.22u 1 2
Rp 1 2 372.838
Cp 1 2 9.315p
Rs 1 N3 0.00037
L1 N3 2 0.214797u
.ends 1010P_7443936050022_0.22u
*******
.subckt 1010P_7443936050068_0.68u 1 2
Rp 1 2 926.896
Cp 1 2 14.804p
Rs 1 N3 0.00077
L1 N3 2 0.686714u
.ends 1010P_7443936050068_0.68u
*******
.subckt 1010P_744393605010_1u 1 2
Rp 1 2 1119
Cp 1 2 17.716p
Rs 1 N3 0.00097
L1 N3 2 1.03u
.ends 1010P_744393605010_1u
*******
.subckt 1010P_744393605015_1.5u 1 2
Rp 1 2 1851
Cp 1 2 19.815p
Rs 1 N3 0.0014
L1 N3 2 1.47u
.ends 1010P_744393605015_1.5u
*******
.subckt 1010P_744393605022_2.2u 1 2
Rp 1 2 1968
Cp 1 2 17.455p
Rs 1 N3 0.0019
L1 N3 2 2.108u
.ends 1010P_744393605022_2.2u
*******
.subckt 1010P_744393605033_3.3u 1 2
Rp 1 2 2782
Cp 1 2 24.393p
Rs 1 N3 0.0027
L1 N3 2 3.043u
.ends 1010P_744393605033_3.3u
*******
.subckt 1010P_744393605047_4.7u 1 2
Rp 1 2 2776
Cp 1 2 23.894p
Rs 1 N3 0.0038
L1 N3 2 4.413u
.ends 1010P_744393605047_4.7u
*******
.subckt 1010P_744393605056_5.6u 1 2
Rp 1 2 4293
Cp 1 2 20.905p
Rs 1 N3 0.005
L1 N3 2 5.669u
.ends 1010P_744393605056_5.6u
*******
.subckt 1010P_744393605068_6.8u 1 2
Rp 1 2 4296
Cp 1 2 25.522p
Rs 1 N3 0.0059
L1 N3 2 6.595u
.ends 1010P_744393605068_6.8u
*******
.subckt 1010P_744393605082_8.2u 1 2
Rp 1 2 5160
Cp 1 2 24.052p
Rs 1 N3 0.0071
L1 N3 2 7.867u
.ends 1010P_744393605082_8.2u
*******
.subckt 1010P_744393605100_10u 1 2
Rp 1 2 6434
Cp 1 2 26.859p
Rs 1 N3 0.0085
L1 N3 2 10.006u
.ends 1010P_744393605100_10u
*******
.subckt 1010P_744393605150_15u 1 2
Rp 1 2 7771
Cp 1 2 25.378p
Rs 1 N3 0.0129
L1 N3 2 15.04u
.ends 1010P_744393605150_15u
*******
.subckt 1010P_744393605220_22u 1 2
Rp 1 2 6827
Cp 1 2 31.171p
Rs 1 N3 0.0187
L1 N3 2 21.974u
.ends 1010P_744393605220_22u
*******
.subckt 1060P_744393665010_1u 1 2
Rp 1 2 1252
Cp 1 2 21.593p
Rs 1 N3 0.0015
L1 N3 2 1.068u
.ends 1060P_744393665010_1u
*******
.subckt 1060P_744393665012_1.2u 1 2
Rp 1 2 1765
Cp 1 2 21.758p
Rs 1 N3 0.0018
L1 N3 2 1.339u
.ends 1060P_744393665012_1.2u
*******
.subckt 1060P_744393665015_1.5u 1 2
Rp 1 2 2186
Cp 1 2 18.19p
Rs 1 N3 0.0021
L1 N3 2 1.601u
.ends 1060P_744393665015_1.5u
*******
.subckt 1060P_744393665022_2.2u 1 2
Rp 1 2 2143
Cp 1 2 21.13p
Rs 1 N3 0.0031
L1 N3 2 2.201u
.ends 1060P_744393665022_2.2u
*******
.subckt 1060P_744393665033_3.3u 1 2
Rp 1 2 2077
Cp 1 2 27.749p
Rs 1 N3 0.0046
L1 N3 2 3.38u
.ends 1060P_744393665033_3.3u
*******
.subckt 1060P_744393665047_4.7u 1 2
Rp 1 2 2945
Cp 1 2 29.968p
Rs 1 N3 0.0057
L1 N3 2 4.446u
.ends 1060P_744393665047_4.7u
*******
.subckt 1060P_744393665056_5.6u 1 2
Rp 1 2 2151
Cp 1 2 33.941p
Rs 1 N3 0.0064
L1 N3 2 6.266u
.ends 1060P_744393665056_5.6u
*******
.subckt 1060P_744393665068_6.8u 1 2
Rp 1 2 2498
Cp 1 2 41.472p
Rs 1 N3 0.0071
L1 N3 2 6.48u
.ends 1060P_744393665068_6.8u
*******
.subckt 1060P_744393665082_8.2u 1 2
Rp 1 2 3685
Cp 1 2 29.508p
Rs 1 N3 0.0107
L1 N3 2 8.102u
.ends 1060P_744393665082_8.2u
*******
.subckt 1060P_744393665100_10u 1 2
Rp 1 2 4059
Cp 1 2 31.132p
Rs 1 N3 0.0126
L1 N3 2 9.703u
.ends 1060P_744393665100_10u
*******
.subckt 1090_74439369010_1u 1 2
Rp 1 2 1136
Cp 1 2 14.279p
Rs 1 N3 0.0014
L1 N3 2 1.069u
.ends 1090_74439369010_1u
*******
.subckt 1090_74439369015_1.5u 1 2
Rp 1 2 1195
Cp 1 2 19.206p
Rs 1 N3 0.00146
L1 N3 2 1.349u
.ends 1090_74439369015_1.5u
*******
.subckt 1090_74439369022_2.2u 1 2
Rp 1 2 2074
Cp 1 2 14.601p
Rs 1 N3 0.0022
L1 N3 2 2.242u
.ends 1090_74439369022_2.2u
*******
.subckt 1090_74439369033_3.3u 1 2
Rp 1 2 3017
Cp 1 2 14.697p
Rs 1 N3 0.0034
L1 N3 2 3.164u
.ends 1090_74439369033_3.3u
*******
.subckt 1090_74439369047_4.7u 1 2
Rp 1 2 4114
Cp 1 2 12.704p
Rs 1 N3 0.005
L1 N3 2 4.625u
.ends 1090_74439369047_4.7u
*******
.subckt 1090_74439369056_5.6u 1 2
Rp 1 2 4898
Cp 1 2 13.52p
Rs 1 N3 0.0059
L1 N3 2 5.491u
.ends 1090_74439369056_5.6u
*******
.subckt 1090_74439369068_6.8u 1 2
Rp 1 2 5791
Cp 1 2 14.891p
Rs 1 N3 0.00716
L1 N3 2 7.08u
.ends 1090_74439369068_6.8u
*******
.subckt 1090_74439369082_8.2u 1 2
Rp 1 2 7214
Cp 1 2 12.059p
Rs 1 N3 0.01
L1 N3 2 8.743u
.ends 1090_74439369082_8.2u
*******
.subckt 1090_74439369100_10u 1 2
Rp 1 2 7876
Cp 1 2 13.203p
Rs 1 N3 0.011
L1 N3 2 10.09u
.ends 1090_74439369100_10u
*******
.subckt 1090_74439369150_15u 1 2
Rp 1 2 8204
Cp 1 2 14.622p
Rs 1 N3 0.0148
L1 N3 2 14.546u
.ends 1090_74439369150_15u
*******
.subckt 1090_74439369220_22u 1 2
Rp 1 2 10223
Cp 1 2 16.595p
Rs 1 N3 0.021
L1 N3 2 20.401u
.ends 1090_74439369220_22u
*******
.subckt 1090_74439369330_33u 1 2
Rp 1 2 9749
Cp 1 2 16.728p
Rs 1 N3 0.0362
L1 N3 2 32.37u
.ends 1090_74439369330_33u
*******
.subckt 1510_74439370033_3.3u 1 2
Rp 1 2 2766
Cp 1 2 30.279p
Rs 1 N3 0.0026
L1 N3 2 3.298u
.ends 1510_74439370033_3.3u
*******
.subckt 1510_74439370047_4.7u 1 2
Rp 1 2 4296
Cp 1 2 22.242p
Rs 1 N3 0.0031
L1 N3 2 4.217u
.ends 1510_74439370047_4.7u
*******
.subckt 1510_74439370056_5.6u 1 2
Rp 1 2 3418
Cp 1 2 30.225p
Rs 1 N3 0.0035
L1 N3 2 5.283u
.ends 1510_74439370056_5.6u
*******
.subckt 1510_74439370068_6.8u 1 2
Rp 1 2 5066
Cp 1 2 21.801p
Rs 1 N3 0.0041
L1 N3 2 6.111u
.ends 1510_74439370068_6.8u
*******
.subckt 1510_74439370082_8.2u 1 2
Rp 1 2 6284
Cp 1 2 25.54p
Rs 1 N3 0.0055
L1 N3 2 8.328u
.ends 1510_74439370082_8.2u
*******
.subckt 1510_74439370100_10u 1 2
Rp 1 2 5244
Cp 1 2 29.045p
Rs 1 N3 0.0064
L1 N3 2 10.4u
.ends 1510_74439370100_10u
*******
.subckt 1510_74439370150_15u 1 2
Rp 1 2 7827
Cp 1 2 24.013p
Rs 1 N3 0.0105
L1 N3 2 15.895u
.ends 1510_74439370150_15u
*******
.subckt 1510_74439370220_22u 1 2
Rp 1 2 8204
Cp 1 2 26.195p
Rs 1 N3 0.0125
L1 N3 2 20.695u
.ends 1510_74439370220_22u
*******
.subckt 1510_74439370330_33u 1 2
Rp 1 2 10776
Cp 1 2 27.127p
Rs 1 N3 0.018
L1 N3 2 31.904u
.ends 1510_74439370330_33u
*******
.subckt 4020_744393230011_0.11u 1 2
Rp 1 2 301
Cp 1 2 2p
Rs 1 N3 0.002
L1 N3 2 0.106u
.ends 4020_744393230011_0.11u
*******
.subckt 4020_744393230022_0.22u 1 2
Rp 1 2 500
Cp 1 2 4.1p
Rs 1 N3 0.00305
L1 N3 2 0.231u
.ends 4020_744393230022_0.22u
*******
.subckt 4020_744393230047_0.47u 1 2
Rp 1 2 560.457
Cp 1 2 5.571p
Rs 1 N3 0.00525
L1 N3 2 0.47u
.ends 4020_744393230047_0.47u
*******
.subckt 4020_744393230056_0.56u 1 2
Rp 1 2 1264
Cp 1 2 6.009p
Rs 1 N3 0.0063
L1 N3 2 0.54u
.ends 4020_744393230056_0.56u
*******
.subckt 4020_744393230068_0.68u 1 2
Rp 1 2 1050
Cp 1 2 6.38p
Rs 1 N3 0.0066
L1 N3 2 0.63u
.ends 4020_744393230068_0.68u
*******
.subckt 4020_744393230082_0.82u 1 2
Rp 1 2 1325
Cp 1 2 6.414p
Rs 1 N3 0.0093
L1 N3 2 0.81u
.ends 4020_744393230082_0.82u
*******
.subckt 4020_74439323010_1u 1 2
Rp 1 2 1442
Cp 1 2 7.529p
Rs 1 N3 0.0107
L1 N3 2 1.03u
.ends 4020_74439323010_1u
*******
.subckt 4020_74439323012_1.2u 1 2
Rp 1 2 1678
Cp 1 2 7.325p
Rs 1 N3 0.0125
L1 N3 2 1.17u
.ends 4020_74439323012_1.2u
*******
.subckt 4020_74439323015_1.5u 1 2
Rp 1 2 2102
Cp 1 2 6.133p
Rs 1 N3 0.0163
L1 N3 2 1.44u
.ends 4020_74439323015_1.5u
*******
.subckt 4020_74439323022_2.2u 1 2
Rp 1 2 3075
Cp 1 2 8.237p
Rs 1 N3 0.0202
L1 N3 2 2.25u
.ends 4020_74439323022_2.2u
*******
.subckt 4030_744393240033_0.33u 1 2
Rp 1 2 457
Cp 1 2 6p
Rs 1 N3 0.0031
L1 N3 2 0.314u
.ends 4030_744393240033_0.33u
*******
.subckt 4030_744393240047_0.47u 1 2
Rp 1 2 707.603
Cp 1 2 5.023p
Rs 1 N3 0.0039
L1 N3 2 0.444u
.ends 4030_744393240047_0.47u
*******
.subckt 4030_744393240056_0.56u 1 2
Rp 1 2 981.099
Cp 1 2 5.572p
Rs 1 N3 0.0041
L1 N3 2 0.59u
.ends 4030_744393240056_0.56u
*******
.subckt 4030_744393240064_0.64u 1 2
Rp 1 2 1004
Cp 1 2 5.533p
Rs 1 N3 0.0048
L1 N3 2 0.591u
.ends 4030_744393240064_0.64u
*******
.subckt 4030_74439324010_1u 1 2
Rp 1 2 1294
Cp 1 2 7.665p
Rs 1 N3 0.0087
L1 N3 2 0.65u
.ends 4030_74439324010_1u
*******
.subckt 4030_744393240090_0.90u 1 2
Rp 1 2 1043
Cp 1 2 7.898p
Rs 1 N3 0.0061
L1 N3 2 0.84u
.ends 4030_744393240090_0.90u
*******
.subckt 4030_74439324012_1.2u 1 2
Rp 1 2 1507
Cp 1 2 7.672p
Rs 1 N3 0.0089
L1 N3 2 1.19u
.ends 4030_74439324012_1.2u
*******
.subckt 4030_74439324015_1.5u 1 2
Rp 1 2 1631
Cp 1 2 6.572p
Rs 1 N3 0.0101
L1 N3 2 1.37u
.ends 4030_74439324015_1.5u
*******
.subckt 4030_74439324022_2.2u 1 2
Rp 1 2 2709
Cp 1 2 7.314p
Rs 1 N3 0.0166
L1 N3 2 2.12u
.ends 4030_74439324022_2.2u
*******
.subckt 4030_74439324033_3.3u 1 2
Rp 1 2 2911
Cp 1 2 8.896p
Rs 1 N3 0.0202
L1 N3 2 3.26u
.ends 4030_74439324033_3.3u
*******
.subckt 4030_74439324047_4.7u 1 2
Rp 1 2 6900
Cp 1 2 7.185p
Rs 1 N3 0.0313
L1 N3 2 4.49u
.ends 4030_74439324047_4.7u
*******
.subckt 4040_74439325033_3.3u 1 2
Rp 1 2 2925
Cp 1 2 8.544p
Rs 1 N3 0.0204
L1 N3 2 3.217u
.ends 4040_74439325033_3.3u
*******
.subckt 4040_74439325047_4.7u 1 2
Rp 1 2 2552
Cp 1 2 9.462p
Rs 1 N3 0.0265
L1 N3 2 4.966u
.ends 4040_74439325047_4.7u
*******
.subckt 4040_74439325056_5.6u 1 2
Rp 1 2 6407
Cp 1 2 8.287p
Rs 1 N3 0.0342
L1 N3 2 5.719u
.ends 4040_74439325056_5.6u
*******
.subckt 4040_74439325068_6.8u 1 2
Rp 1 2 10604
Cp 1 2 6.978p
Rs 1 N3 0.0423
L1 N3 2 6.707u
.ends 4040_74439325068_6.8u
*******
.subckt 5020_744393330016_0.16u 1 2
Rp 1 2 332.836
Cp 1 2 4.771p
Rs 1 N3 0.0022
L1 N3 2 0.148u
.ends 5020_744393330016_0.16u
*******
.subckt 5020_744393330033_0.33u 1 2
Rp 1 2 546.947
Cp 1 2 7.165p
Rs 1 N3 0.003
L1 N3 2 0.332u
.ends 5020_744393330033_0.33u
*******
.subckt 5020_744393330056_0.56u 1 2
Rp 1 2 849.046
Cp 1 2 5.993p
Rs 1 N3 0.0052
L1 N3 2 0.536u
.ends 5020_744393330056_0.56u
*******
.subckt 5020_744393330068_0.68u 1 2
Rp 1 2 1181
Cp 1 2 6.54p
Rs 1 N3 0.0067
L1 N3 2 0.72u
.ends 5020_744393330068_0.68u
*******
.subckt 5020_74439333010_1u 1 2
Rp 1 2 950
Cp 1 2 9.636p
Rs 1 N3 0.0095
L1 N3 2 0.97u
.ends 5020_74439333010_1u
*******
.subckt 5020_74439333012_1.2u 1 2
Rp 1 2 1708
Cp 1 2 8.409p
Rs 1 N3 0.0108
L1 N3 2 1.25u
.ends 5020_74439333012_1.2u
*******
.subckt 5030_744393340016_0.16u 1 2
Rp 1 2 335
Cp 1 2 4.509p
Rs 1 N3 0.0021
L1 N3 2 0.154u
.ends 5030_744393340016_0.16u
*******
.subckt 5030_744393340033_0.33u 1 2
Rp 1 2 574.378
Cp 1 2 7.026p
Rs 1 N3 0.00301
L1 N3 2 0.328238u
.ends 5030_744393340033_0.33u
*******
.subckt 5030_744393340056_0.56u 1 2
Rp 1 2 836.509
Cp 1 2 8.126p
Rs 1 N3 0.00399
L1 N3 2 0.546969u
.ends 5030_744393340056_0.56u
*******
.subckt 5030_74439334010_1u 1 2
Rp 1 2 810.15
Cp 1 2 10.541p
Rs 1 N3 0.0063
L1 N3 2 0.66854u
.ends 5030_74439334010_1u
*******
.subckt 5030_744393340068_0.68u 1 2
Rp 1 2 613.431
Cp 1 2 9.363p
Rs 1 N3 0.00409
L1 N3 2 0.691759u
.ends 5030_744393340068_0.68u
*******
.subckt 5030_74439334012_1.2u 1 2
Rp 1 2 1486
Cp 1 2 9.582p
Rs 1 N3 0.0066
L1 N3 2 1.219u
.ends 5030_74439334012_1.2u
*******
.subckt 5030_74439334015_1.5u 1 2
Rp 1 2 1932
Cp 1 2 8.871p
Rs 1 N3 0.008
L1 N3 2 1.614u
.ends 5030_74439334015_1.5u
*******
.subckt 5030_74439334018_1.8u 1 2
Rp 1 2 2463
Cp 1 2 8.913p
Rs 1 N3 0.0091
L1 N3 2 1.88u
.ends 5030_74439334018_1.8u
*******
.subckt 5030_74439334022_2.2u 1 2
Rp 1 2 2762
Cp 1 2 9.83p
Rs 1 N3 0.0113
L1 N3 2 2.13u
.ends 5030_74439334022_2.2u
*******
.subckt 5030_74439334033_3.3u 1 2
Rp 1 2 2140
Cp 1 2 11.045p
Rs 1 N3 0.0163
L1 N3 2 3.496u
.ends 5030_74439334033_3.3u
*******
.subckt 5030_74439334047_4.7u 1 2
Rp 1 2 3991
Cp 1 2 10.549p
Rs 1 N3 0.0229
L1 N3 2 4.943u
.ends 5030_74439334047_4.7u
*******
.subckt 5050_744393305033_3.3u 1 2
Rp 1 2 1606
Cp 1 2 11.453p
Rs 1 N3 0.0132
L1 N3 2 3.213u
.ends 5050_744393305033_3.3u
*******
.subckt 5050_744393305056_5.6u 1 2
Rp 1 2 3527
Cp 1 2 9.72p
Rs 1 N3 0.0218
L1 N3 2 5.702u
.ends 5050_744393305056_5.6u
*******
.subckt 5050_744393305068_6.8u 1 2
Rp 1 2 9422
Cp 1 2 11.47p
Rs 1 N3 0.0237
L1 N3 2 6.846u
.ends 5050_744393305068_6.8u
*******
.subckt 5050_744393305082_8.2u 1 2
Rp 1 2 11476
Cp 1 2 10.965p
Rs 1 N3 0.0293
L1 N3 2 8.338u
.ends 5050_744393305082_8.2u
*******
.subckt 5050_744393305100_10u 1 2
Rp 1 2 4502
Cp 1 2 12.201p
Rs 1 N3 0.0354
L1 N3 2 10.647u
.ends 5050_744393305100_10u
*******
.subckt 5050_744393305150_15u 1 2
Rp 1 2 17051
Cp 1 2 10.749p
Rs 1 N3 0.0568
L1 N3 2 16.504u
.ends 5050_744393305150_15u
*******
.subckt 5050_744393305220_22u 1 2
Rp 1 2 19323
Cp 1 2 11.699p
Rs 1 N3 0.075
L1 N3 2 22.094u
.ends 5050_744393305220_22u
*******
.subckt 6030_744393440015_0.15u 1 2
Rp 1 2 306.09
Cp 1 2 4.722p
Rs 1 N3 0.00124
L1 N3 2 0.147u
.ends 6030_744393440015_0.15u
*******
.subckt 6030_744393440018_0.18u 1 2
Rp 1 2 393.041
Cp 1 2 5.062p
Rs 1 N3 0.00132
L1 N3 2 0.176u
.ends 6030_744393440018_0.18u
*******
.subckt 6030_744393440033_0.33u 1 2
Rp 1 2 683.781
Cp 1 2 6.324p
Rs 1 N3 0.0021
L1 N3 2 0.316u
.ends 6030_744393440033_0.33u
*******
.subckt 6030_744393440047_0.47u 1 2
Rp 1 2 708
Cp 1 2 7.228p
Rs 1 N3 0.0028
L1 N3 2 0.469u
.ends 6030_744393440047_0.47u
*******
.subckt 6030_744393440056_0.56u 1 2
Rp 1 2 876.79
Cp 1 2 7.515p
Rs 1 N3 0.0029
L1 N3 2 0.561u
.ends 6030_744393440056_0.56u
*******
.subckt 6030_744393440068_0.68u 1 2
Rp 1 2 853
Cp 1 2 8.355p
Rs 1 N3 0.0038
L1 N3 2 0.713u
.ends 6030_744393440068_0.68u
*******
.subckt 6030_74439344010_1u 1 2
Rp 1 2 1956
Cp 1 2 7.102p
Rs 1 N3 0.0055
L1 N3 2 1.008u
.ends 6030_74439344010_1u
*******
.subckt 6030_74439344012_1.2u 1 2
Rp 1 2 2178
Cp 1 2 8.182p
Rs 1 N3 0.0064
L1 N3 2 1.105u
.ends 6030_74439344012_1.2u
*******
.subckt 6030_74439344018_1.8u 1 2
Rp 1 2 2033
Cp 1 2 8.954p
Rs 1 N3 0.0097
L1 N3 2 1.872u
.ends 6030_74439344018_1.8u
*******
.subckt 6030_74439344022_2.2u 1 2
Rp 1 2 2927
Cp 1 2 8.36p
Rs 1 N3 0.0105
L1 N3 2 2.182u
.ends 6030_74439344022_2.2u
*******
.subckt 6030_74439344033_3.3u 1 2
Rp 1 2 4970
Cp 1 2 7.979p
Rs 1 N3 0.0192
L1 N3 2 3.247u
.ends 6030_74439344033_3.3u
*******
.subckt 6030_74439344047_4.7u 1 2
Rp 1 2 7211
Cp 1 2 7.002p
Rs 1 N3 0.031
L1 N3 2 4.676u
.ends 6030_74439344047_4.7u
*******
.subckt 6030P_7443934450015_0.15u 1 2
Rp 1 2 281.192
Cp 1 2 6.38p
Rs 1 N3 0.0009
L1 N3 2 0.158317u
.ends 6030P_7443934450015_0.15u
*******
.subckt 6030P_7443934450022_0.22u 1 2
Rp 1 2 268.007
Cp 1 2 8.214p
Rs 1 N3 0.0012
L1 N3 2 0.202144u
.ends 6030P_7443934450022_0.22u
*******
.subckt 6030P_7443934450033_0.33u 1 2
Rp 1 2 455.475
Cp 1 2 9.03p
Rs 1 N3 0.0016
L1 N3 2 0.349571u
.ends 6030P_7443934450033_0.33u
*******
.subckt 6030P_7443934450047_0.47u 1 2
Rp 1 2 729.668
Cp 1 2 9.466p
Rs 1 N3 0.0021
L1 N3 2 0.473657u
.ends 6030P_7443934450047_0.47u
*******
.subckt 6030P_7443934450056_0.56u 1 2
Rp 1 2 929.081
Cp 1 2 9.847p
Rs 1 N3 0.0027
L1 N3 2 0.57528u
.ends 6030P_7443934450056_0.56u
*******
.subckt 6030P_7443934450068_0.68u 1 2
Rp 1 2 793.567
Cp 1 2 11.486p
Rs 1 N3 0.0028
L1 N3 2 0.70047u
.ends 6030P_7443934450068_0.68u
*******
.subckt 6030P_7443934450082_0.82u 1 2
Rp 1 2 978.457
Cp 1 2 12.258p
Rs 1 N3 0.0034
L1 N3 2 0.829331u
.ends 6030P_7443934450082_0.82u
*******
.subckt 6030P_744393445010_1u 1 2
Rp 1 2 1160
Cp 1 2 9.957p
Rs 1 N3 0.0042
L1 N3 2 1.021u
.ends 6030P_744393445010_1u
*******
.subckt 6030P_744393445012_1.2u 1 2
Rp 1 2 1132
Cp 1 2 11.176p
Rs 1 N3 0.0043
L1 N3 2 1.149u
.ends 6030P_744393445012_1.2u
*******
.subckt 6030P_744393445015_1.5u 1 2
Rp 1 2 1939
Cp 1 2 16.6p
Rs 1 N3 0.0058
L1 N3 2 1.389u
.ends 6030P_744393445015_1.5u
*******
.subckt 6030P_744393445018_1.8u 1 2
Rp 1 2 1665
Cp 1 2 17.179p
Rs 1 N3 0.0068
L1 N3 2 1.906u
.ends 6030P_744393445018_1.8u
*******
.subckt 6030P_744393445022_2.2u 1 2
Rp 1 2 2086
Cp 1 2 14.921p
Rs 1 N3 0.0083
L1 N3 2 2.194u
.ends 6030P_744393445022_2.2u
*******
.subckt 6030P_744393445033_3.3u 1 2
Rp 1 2 2368
Cp 1 2 15.869p
Rs 1 N3 0.0143
L1 N3 2 3.294u
.ends 6030P_744393445033_3.3u
*******
.subckt 6030P_744393445047_4.7u 1 2
Rp 1 2 3260
Cp 1 2 17.613p
Rs 1 N3 0.0167
L1 N3 2 4.738u
.ends 6030P_744393445047_4.7u
*******
.subckt 6030P_744393445056_5.6u 1 2
Rp 1 2 1705
Cp 1 2 21.665p
Rs 1 N3 0.0199
L1 N3 2 4.867u
.ends 6030P_744393445056_5.6u
*******
.subckt 6030P_744393445068_6.8u 1 2
Rp 1 2 3986
Cp 1 2 17.868p
Rs 1 N3 0.0244
L1 N3 2 5.901u
.ends 6030P_744393445068_6.8u
*******
.subckt 6030P_744393445082_8.2u 1 2
Rp 1 2 5343
Cp 1 2 14.909p
Rs 1 N3 0.036
L1 N3 2 7.949u
.ends 6030P_744393445082_8.2u
*******
.subckt 6030P_744393445100_10u 1 2
Rp 1 2 5158
Cp 1 2 15.729p
Rs 1 N3 0.0403
L1 N3 2 9.521u
.ends 6030P_744393445100_10u
*******
.subckt 6030P_744393445120_12u 1 2
Rp 1 2 5255
Cp 1 2 16.483p
Rs 1 N3 0.0485
L1 N3 2 11.479u
.ends 6030P_744393445120_12u
*******
.subckt 6030P_744393445150_15u 1 2
Rp 1 2 5431
Cp 1 2 21.205p
Rs 1 N3 0.0618
L1 N3 2 16.013u
.ends 6030P_744393445150_15u
*******
.subckt 6030P_744393445180_18u 1 2
Rp 1 2 5251
Cp 1 2 22.753p
Rs 1 N3 0.0683
L1 N3 2 18.856u
.ends 6030P_744393445180_18u
*******
.subckt 6060_74439346010_1u 1 2
Rp 1 2 1210
Cp 1 2 6.845p
Rs 1 N3 0.00339
L1 N3 2 1.046u
.ends 6060_74439346010_1u
*******
.subckt 6060_74439346012_1.2u 1 2
Rp 1 2 1330
Cp 1 2 8.78p
Rs 1 N3 0.00365
L1 N3 2 1.158u
.ends 6060_74439346012_1.2u
*******
.subckt 6060_74439346015_1.5u 1 2
Rp 1 2 1396
Cp 1 2 9.359p
Rs 1 N3 0.0039
L1 N3 2 1.373u
.ends 6060_74439346015_1.5u
*******
.subckt 6060_74439346018_1.8u 1 2
Rp 1 2 1659
Cp 1 2 7.994p
Rs 1 N3 0.0047
L1 N3 2 1.806u
.ends 6060_74439346018_1.8u
*******
.subckt 6060_74439346022_2.2u 1 2
Rp 1 2 1877
Cp 1 2 8.362p
Rs 1 N3 0.00558
L1 N3 2 2.182u
.ends 6060_74439346022_2.2u
*******
.subckt 6060_74439346033_3.3u 1 2
Rp 1 2 2955
Cp 1 2 8.785p
Rs 1 N3 0.01083
L1 N3 2 2.95u
.ends 6060_74439346033_3.3u
*******
.subckt 6060_74439346047_4.7u 1 2
Rp 1 2 4305
Cp 1 2 7.633p
Rs 1 N3 0.013
L1 N3 2 4.289u
.ends 6060_74439346047_4.7u
*******
.subckt 6060_74439346056_5.6u 1 2
Rp 1 2 5112
Cp 1 2 7.79p
Rs 1 N3 0.015
L1 N3 2 5.311u
.ends 6060_74439346056_5.6u
*******
.subckt 6060_74439346068_6.8u 1 2
Rp 1 2 5867
Cp 1 2 7.976p
Rs 1 N3 0.0176
L1 N3 2 6.553u
.ends 6060_74439346068_6.8u
*******
.subckt 6060_74439346082_8.2u 1 2
Rp 1 2 6820
Cp 1 2 8.668p
Rs 1 N3 0.023
L1 N3 2 7.855u
.ends 6060_74439346082_8.2u
*******
.subckt 6060_74439346100_10u 1 2
Rp 1 2 9786
Cp 1 2 8.192p
Rs 1 N3 0.0265
L1 N3 2 9.539u
.ends 6060_74439346100_10u
*******
.subckt 6060_74439346150_15u 1 2
Rp 1 2 11178
Cp 1 2 8.829p
Rs 1 N3 0.042
L1 N3 2 15.089u
.ends 6060_74439346150_15u
*******
.subckt 6060P_7443934650022_0.22u 1 2
Rp 1 2 684.147
Cp 1 2 7.285p
Rs 1 N3 0.0011
L1 N3 2 0.227919u
.ends 6060P_7443934650022_0.22u
*******
.subckt 6060P_7443934650047_0.47u 1 2
Rp 1 2 602.157
Cp 1 2 8.922p
Rs 1 N3 0.0014
L1 N3 2 0.502539u
.ends 6060P_7443934650047_0.47u
*******
.subckt 6060P_7443934650068_0.68u 1 2
Rp 1 2 608.07
Cp 1 2 9.93p
Rs 1 N3 0.0017
L1 N3 2 0.641243u
.ends 6060P_7443934650068_0.68u
*******
.subckt 6060P_744393465010_1u 1 2
Rp 1 2 900.677
Cp 1 2 12.235p
Rs 1 N3 0.0022
L1 N3 2 1.05u
.ends 6060P_744393465010_1u
*******
.subckt 6060P_744393465012_1.2u 1 2
Rp 1 2 1119
Cp 1 2 14.265p
Rs 1 N3 0.0026
L1 N3 2 1.279u
.ends 6060P_744393465012_1.2u
*******
.subckt 6060P_744393465015_1.5u 1 2
Rp 1 2 891.855
Cp 1 2 17.044p
Rs 1 N3 0.003
L1 N3 2 1.52u
.ends 6060P_744393465015_1.5u
*******
.subckt 6060P_744393465018_1.8u 1 2
Rp 1 2 1198
Cp 1 2 14.596p
Rs 1 N3 0.0035
L1 N3 2 1.775u
.ends 6060P_744393465018_1.8u
*******
.subckt 6060P_744393465022_2.2u 1 2
Rp 1 2 1177
Cp 1 2 12.743p
Rs 1 N3 0.0039
L1 N3 2 2.286u
.ends 6060P_744393465022_2.2u
*******
.subckt 6060P_744393465033_3.3u 1 2
Rp 1 2 1544
Cp 1 2 17.52p
Rs 1 N3 0.006
L1 N3 2 3.353u
.ends 6060P_744393465033_3.3u
*******
.subckt 6060P_744393465047_4.7u 1 2
Rp 1 2 2269
Cp 1 2 13.11p
Rs 1 N3 0.0094
L1 N3 2 4.481u
.ends 6060P_744393465047_4.7u
*******
.subckt 6060P_744393465056_5.6u 1 2
Rp 1 2 2589
Cp 1 2 18.351p
Rs 1 N3 0.0109
L1 N3 2 5.746u
.ends 6060P_744393465056_5.6u
*******
.subckt 6060P_744393465068_6.8u 1 2
Rp 1 2 1882
Cp 1 2 22.539p
Rs 1 N3 0.0125
L1 N3 2 6.644u
.ends 6060P_744393465068_6.8u
*******
.subckt 6060P_744393465082_8.2u 1 2
Rp 1 2 2401
Cp 1 2 20.981p
Rs 1 N3 0.0146
L1 N3 2 8.023u
.ends 6060P_744393465082_8.2u
*******
.subckt 6060P_744393465100_10u 1 2
Rp 1 2 3239
Cp 1 2 18.492p
Rs 1 N3 0.018
L1 N3 2 9.103u
.ends 6060P_744393465100_10u
*******
.subckt 6060P_744393465120_12u 1 2
Rp 1 2 4738
Cp 1 2 16.735p
Rs 1 N3 0.0228
L1 N3 2 11.306u
.ends 6060P_744393465120_12u
*******
.subckt 6060P_744393465150_15u 1 2
Rp 1 2 2569
Cp 1 2 26.54p
Rs 1 N3 0.0286
L1 N3 2 14.381u
.ends 6060P_744393465150_15u
*******
.subckt 6060P_744393465180_18u 1 2
Rp 1 2 2428
Cp 1 2 28.695p
Rs 1 N3 0.0345
L1 N3 2 16.806u
.ends 6060P_744393465180_18u
*******
.subckt 6060P_744393465220_22u 1 2
Rp 1 2 3755
Cp 1 2 18.501p
Rs 1 N3 0.042
L1 N3 2 20.631u
.ends 6060P_744393465220_22u
*******
.subckt 7030_74439384010_1u 1 2
Rp 1 2 1583
Cp 1 2 11.684p
Rs 1 N3 0.0039
L1 N3 2 0.9456u
.ends 7030_74439384010_1u
*******
.subckt 7030_74439384012_1.2u 1 2
Rp 1 2 841
Cp 1 2 14.189p
Rs 1 N3 0.0042
L1 N3 2 1.157u
.ends 7030_74439384012_1.2u
*******
.subckt 7030_74439384015_1.5u 1 2
Rp 1 2 1847
Cp 1 2 11.892p
Rs 1 N3 0.0051
L1 N3 2 1.393u
.ends 7030_74439384015_1.5u
*******
.subckt 7030_74439384022_2.2u 1 2
Rp 1 2 2530
Cp 1 2 14.021p
Rs 1 N3 0.0079
L1 N3 2 2.223u
.ends 7030_74439384022_2.2u
*******
.subckt 7030_74439384033_3.3u 1 2
Rp 1 2 3242
Cp 1 2 12.561p
Rs 1 N3 0.0144
L1 N3 2 3.171u
.ends 7030_74439384033_3.3u
*******
.subckt 7030_74439384047_4.7u 1 2
Rp 1 2 5033
Cp 1 2 13.362p
Rs 1 N3 0.0198
L1 N3 2 5.149u
.ends 7030_74439384047_4.7u
*******
.subckt 7070_74439387033_3.3u 1 2
Rp 1 2 2426
Cp 1 2 14.688p
Rs 1 N3 0.0064
L1 N3 2 3.212u
.ends 7070_74439387033_3.3u
*******
.subckt 7070_74439387047_4.7u 1 2
Rp 1 2 3245
Cp 1 2 13.478p
Rs 1 N3 0.0092
L1 N3 2 4.617u
.ends 7070_74439387047_4.7u
*******
.subckt 7070_74439387056_5.6u 1 2
Rp 1 2 2248
Cp 1 2 18.924p
Rs 1 N3 0.0124
L1 N3 2 5.67u
.ends 7070_74439387056_5.6u
*******
.subckt 7070_74439387068_6.8u 1 2
Rp 1 2 2887
Cp 1 2 15.001p
Rs 1 N3 0.0124
L1 N3 2 6.749u
.ends 7070_74439387068_6.8u
*******
.subckt 7070_74439387082_8.2u 1 2
Rp 1 2 3645
Cp 1 2 16.219p
Rs 1 N3 0.0145
L1 N3 2 8.537u
.ends 7070_74439387082_8.2u
*******
.subckt 7070_74439387100_10u 1 2
Rp 1 2 4865
Cp 1 2 14.504p
Rs 1 N3 0.019
L1 N3 2 9.866u
.ends 7070_74439387100_10u
*******
.subckt 8080_744393580068_0.68u 1 2
Rp 1 2 1027
Cp 1 2 9.182p
Rs 1 N3 0.00141
L1 N3 2 0.71u
.ends 8080_744393580068_0.68u
*******
.subckt 8080_74439358010_1u 1 2
Rp 1 2 1445
Cp 1 2 8.916p
Rs 1 N3 0.0021
L1 N3 2 1.014u
.ends 8080_74439358010_1u
*******
.subckt 8080_74439358015_1.5u 1 2
Rp 1 2 1599
Cp 1 2 11.49p
Rs 1 N3 0.00291
L1 N3 2 1.588u
.ends 8080_74439358015_1.5u
*******
.subckt 8080_74439358022_2.2u 1 2
Rp 1 2 2282
Cp 1 2 10.434p
Rs 1 N3 0.0037
L1 N3 2 2.209u
.ends 8080_74439358022_2.2u
*******
.subckt 8080_74439358033_3.3u 1 2
Rp 1 2 2961
Cp 1 2 10.892p
Rs 1 N3 0.0068
L1 N3 2 3.584u
.ends 8080_74439358033_3.3u
*******
.subckt 8080_74439358047_4.7u 1 2
Rp 1 2 4439
Cp 1 2 10.924p
Rs 1 N3 0.00865
L1 N3 2 4.785u
.ends 8080_74439358047_4.7u
*******
.subckt 8080_74439358068_6.8u 1 2
Rp 1 2 6545
Cp 1 2 7.924p
Rs 1 N3 0.013
L1 N3 2 6.596u
.ends 8080_74439358068_6.8u
*******
.subckt 8080_74439358100_10u 1 2
Rp 1 2 8417
Cp 1 2 8.116p
Rs 1 N3 0.019
L1 N3 2 10.282u
.ends 8080_74439358100_10u
*******
.subckt 8080_74439358150_15u 1 2
Rp 1 2 8485
Cp 1 2 11.885p
Rs 1 N3 0.025
L1 N3 2 14.163u
.ends 8080_74439358150_15u
*******
.subckt 8080_74439358220_22u 1 2
Rp 1 2 6467
Cp 1 2 16.367p
Rs 1 N3 0.0307
L1 N3 2 20.685u
.ends 8080_74439358220_22u
*******
