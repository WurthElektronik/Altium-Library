**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  MLCCs - Multilayer Ceramic Chip Capacitors
* Matchcode:              WCAP-CSGP_6-3V
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/19/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0201_885012004003_1.5pF 1 2
Rser 1 3 0.8126
Lser 2 4 0.00000000022
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0201_885012004003_1.5pF
*******
.subckt 0201_885012004004_10pF 1 2
Rser 1 3 0.6361
Lser 2 4 0.00000000022
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0201_885012004004_10pF
*******
.subckt 0201_885012004005_12pF 1 2
Rser 1 3 0.4731
Lser 2 4 0.00000000021
C1 3 4 0.000000000012
Rpar 3 4 10000000000
.ends 0201_885012004005_12pF
*******
.subckt 0201_885012004006_15pF 1 2
Rser 1 3 0.4471
Lser 2 4 0.00000000025
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0201_885012004006_15pF
*******
.subckt 0201_885012004007_18pF 1 2
Rser 1 3 0.4894
Lser 2 4 0.000000000295
C1 3 4 0.000000000018
Rpar 3 4 10000000000
.ends 0201_885012004007_18pF
*******
.subckt 0201_885012004008_22pF 1 2
Rser 1 3 0.5288
Lser 2 4 0.00000000026
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0201_885012004008_22pF
*******
.subckt 0201_885012004009_33pF 1 2
Rser 1 3 0.3381
Lser 2 4 0.000000000257
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0201_885012004009_33pF
*******
.subckt 0201_885012004010_47pF 1 2
Rser 1 3 0.241
Lser 2 4 0.0000000002
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0201_885012004010_47pF
*******
.subckt 0201_885012004001_100pF 1 2
Rser 1 3 0.2125
Lser 2 4 0.00000000025
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0201_885012004001_100pF
*******
.subckt 0201_885012204006_1nF 1 2
Rser 1 3 0.2367
Lser 2 4 0.000000000173
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0201_885012204006_1nF
*******
.subckt 0201_885012104008_4.7nF 1 2
Rser 1 3 0.093
Lser 2 4 0.000000000212
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0201_885012104008_4.7nF
*******
.subckt 0201_885012204004_10nF 1 2
Rser 1 3 0.0709
Lser 2 4 0.00000000018
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012204004_10nF
*******
.subckt 0201_885012104014_10nF 1 2
Rser 1 3 0.0639
Lser 2 4 0.00000000021
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0201_885012104014_10nF
*******
.subckt 0201_885012104005_100nF 1 2
Rser 1 3 0.0287
Lser 2 4 0.00000000015
C1 3 4 0.0000001
Rpar 3 4 500000000
.ends 0201_885012104005_100nF
*******
.subckt 0402_885012005034_1pF 1 2
Rser 1 3 0.734
Lser 2 4 0.00000000038
C1 3 4 0.000000000001
Rpar 3 4 10000000000
.ends 0402_885012005034_1pF
*******
.subckt 0402_885012005035_1.5pF 1 2
Rser 1 3 0.75
Lser 2 4 0.00000000031
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0402_885012005035_1.5pF
*******
.subckt 0402_885012005037_3.3pF 1 2
Rser 1 3 1.5
Lser 2 4 0.00000000039
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0402_885012005037_3.3pF
*******
.subckt 0402_885012005038_4.7pF 1 2
Rser 1 3 0.46
Lser 2 4 0.000000000365
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0402_885012005038_4.7pF
*******
.subckt 0402_885012005039_6.8pF 1 2
Rser 1 3 0.465
Lser 2 4 0.00000000031
C1 3 4 0.00000000000682
Rpar 3 4 10000000000
.ends 0402_885012005039_6.8pF
*******
.subckt 0402_885012005040_10pF 1 2
Rser 1 3 0.467848447943
Lser 2 4 3.77046381E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005040_10pF
*******
.subckt 0402_885012005041_15pF 1 2
Rser 1 3 0.34552139712
Lser 2 4 3.31461104E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885012005041_15pF
*******
.subckt 0402_885012005042_22pF 1 2
Rser 1 3 0.285282706764
Lser 2 4 3.08207076E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885012005042_22pF
*******
.subckt 0402_885012005043_33pF 1 2
Rser 1 3 0.230231956882
Lser 2 4 2.96875149E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005043_33pF
*******
.subckt 0402_885012005044_47pF 1 2
Rser 1 3 0.203455175683
Lser 2 4 3.46537476E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005044_47pF
*******
.subckt 0402_885012005045_68pF 1 2
Rser 1 3 0.18781473697
Lser 2 4 3.22027908E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005045_68pF
*******
.subckt 0402_885012005046_100pF 1 2
Rser 1 3 0.0759217345208
Lser 2 4 3.94922966E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005046_100pF
*******
.subckt 0402_885012005047_150pF 1 2
Rser 1 3 0.112246046138
Lser 2 4 2.15549473E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012005047_150pF
*******
.subckt 0402_885012005048_220pF 1 2
Rser 1 3 0.104232515193
Lser 2 4 1.92172989E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012005048_220pF
*******
.subckt 0402_885012105018_100nF 1 2
Rser 1 3 0.026120802334
Lser 2 4 3.09671131E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012105018_100nF
*******
.subckt 0402_885012205038_100pF 1 2
Rser 1 3 0.81685
Lser 2 4 0.00000000015556
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012205038_100pF
*******
.subckt 0402_885012205039_150pF 1 2
Rser 1 3 0.63099
Lser 2 4 0.00000000012911
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012205039_150pF
*******
.subckt 0402_885012205040_220pF 1 2
Rser 1 3 0.56531
Lser 2 4 0.00000000019063
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012205040_220pF
*******
.subckt 0402_885012205041_330pF 1 2
Rser 1 3 0.47337
Lser 2 4 0.00000000018072
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012205041_330pF
*******
.subckt 0402_885012205042_470pF 1 2
Rser 1 3 0.34662
Lser 2 4 0.00000000017045
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012205042_470pF
*******
.subckt 0402_885012205043_680pF 1 2
Rser 1 3 0.26546
Lser 2 4 0.00000000014081
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0402_885012205043_680pF
*******
.subckt 0402_885012205044_1nF 1 2
Rser 1 3 0.2145
Lser 2 4 0.000000000153
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205044_1nF
*******
.subckt 0402_885012205045_1.5nF 1 2
Rser 1 3 0.20285
Lser 2 4 0.00000000025723
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0402_885012205045_1.5nF
*******
.subckt 0402_885012205046_2.2nF 1 2
Rser 1 3 0.16081
Lser 2 4 0.00000000018799
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0402_885012205046_2.2nF
*******
.subckt 0402_885012205047_3.3nF 1 2
Rser 1 3 0.12518
Lser 2 4 0.00000000020592
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0402_885012205047_3.3nF
*******
.subckt 0402_885012205048_4.7nF 1 2
Rser 1 3 0.09048
Lser 2 4 0.00000000014994
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205048_4.7nF
*******
.subckt 0402_885012205049_6.8nF 1 2
Rser 1 3 0.071
Lser 2 4 0.00000000019016
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0402_885012205049_6.8nF
*******
.subckt 0402_885012205050_10nF 1 2
Rser 1 3 0.0592
Lser 2 4 0.00000000014515
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0402_885012205050_10nF
*******
.subckt 0402_885012205051_15nF 1 2
Rser 1 3 0.03784
Lser 2 4 0.00000000020335
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0402_885012205051_15nF
*******
.subckt 0402_885012205052_22nF 1 2
Rser 1 3 0.0548
Lser 2 4 0.00000000019383
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0402_885012205052_22nF
*******
.subckt 0402_885012205053_33nF 1 2
Rser 1 3 0.03148
Lser 2 4 0.0000000002517
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0402_885012205053_33nF
*******
.subckt 0402_885012205054_47nF 1 2
Rser 1 3 0.02098
Lser 2 4 0.00000000019891
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0402_885012205054_47nF
*******
.subckt 0402_885012205085_100nF 1 2
Rser 1 3 0.035
Lser 2 4 7.65573672E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205085_100nF
*******
.subckt 0402_885012205085R_100nF 1 2
Rser 1 3 0.035
Lser 2 4 7.65573672E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0402_885012205085R_100nF
*******
.subckt 0603_885012006030_4.7pF 1 2
Rser 1 3 0.29124727578
Lser 2 4 4.29705418E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0603_885012006030_4.7pF
*******
.subckt 0603_885012006031_6.8pF 1 2
Rser 1 3 0.299024437013
Lser 2 4 4.5809474E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0603_885012006031_6.8pF
*******
.subckt 0603_885012006032_10pF 1 2
Rser 1 3 0.445774201336
Lser 2 4 4.28073844E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006032_10pF
*******
.subckt 0603_885012006033_15pF 1 2
Rser 1 3 0.353119905486
Lser 2 4 4.35266975E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006033_15pF
*******
.subckt 0603_885012006034_22pF 1 2
Rser 1 3 0.352481322316
Lser 2 4 5.8820344E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006034_22pF
*******
.subckt 0603_885012006035_33pF 1 2
Rser 1 3 0.305919966941
Lser 2 4 5.25713034E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006035_33pF
*******
.subckt 0603_885012006036_47pF 1 2
Rser 1 3 0.062255914612
Lser 2 4 4.24328623E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006036_47pF
*******
.subckt 0603_885012006037_68pF 1 2
Rser 1 3 0.159672910297
Lser 2 4 6.46220787E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006037_68pF
*******
.subckt 0603_885012006038_100pF 1 2
Rser 1 3 0.130130495234
Lser 2 4 5.8979323E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006038_100pF
*******
.subckt 0603_885012006039_150pF 1 2
Rser 1 3 0.097154893647
Lser 2 4 5.82598828E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006039_150pF
*******
.subckt 0603_885012006040_220pF 1 2
Rser 1 3 0.111748485631
Lser 2 4 6.02628009E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012006040_220pF
*******
.subckt 0603_885012006041_330pF 1 2
Rser 1 3 0.0829140919635
Lser 2 4 3.85173897E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006041_330pF
*******
.subckt 0603_885012006042_470pF 1 2
Rser 1 3 0.0647178553788
Lser 2 4 3.67931779E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006042_470pF
*******
.subckt 0603_885012006043_680pF 1 2
Rser 1 3 0.0641029132415
Lser 2 4 3.05763584E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006043_680pF
*******
.subckt 0603_885012006044_1nF 1 2
Rser 1 3 0.0419451701409
Lser 2 4 4.48170961E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006044_1nF
*******
.subckt 0603_885012106019_220nF 1 2
Rser 1 3 0.0108961182185
Lser 2 4 2.50789051E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012106019_220nF
*******
.subckt 0603_885012106020_470nF 1 2
Rser 1 3 0.00976845934589
Lser 2 4 2.50682976E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012106020_470nF
*******
.subckt 0603_885012106021_680nF 1 2
Rser 1 3 0.00991319698945
Lser 2 4 3.55175418E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0603_885012106021_680nF
*******
.subckt 0603_885012106022_1uF 1 2
Rser 1 3 0.00857861035867
Lser 2 4 3.03497279E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0603_885012106022_1uF
*******
.subckt 0603_885012106030_1uF 1 2
Rser 1 3 0.013
Lser 2 4 0.0000000008
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0603_885012106030_1uF
*******
.subckt 0603_885012106031_10uF 1 2
Rser 1 3 0.0105
Lser 2 4 0.0000000008
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 0603_885012106031_10uF
*******
.subckt 0603_885012206053_100pF 1 2
Rser 1 3 0.91003
Lser 2 4 0.00000000024509
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206053_100pF
*******
.subckt 0603_885012206054_150pF 1 2
Rser 1 3 0.68385
Lser 2 4 0.00000000029018
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012206054_150pF
*******
.subckt 0603_885012206055_220pF 1 2
Rser 1 3 0.58631
Lser 2 4 0.00000000033037
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012206055_220pF
*******
.subckt 0603_885012206056_330pF 1 2
Rser 1 3 0.42401
Lser 2 4 0.00000000033129
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206056_330pF
*******
.subckt 0603_885012206057_470pF 1 2
Rser 1 3 0.34594
Lser 2 4 0.00000000033084
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206057_470pF
*******
.subckt 0603_885012206058_680pF 1 2
Rser 1 3 0.29796
Lser 2 4 0.00000000037378
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206058_680pF
*******
.subckt 0603_885012206059_1nF 1 2
Rser 1 3 0.22136
Lser 2 4 0.00000000036253
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206059_1nF
*******
.subckt 0603_885012206060_1.5nF 1 2
Rser 1 3 0.18842
Lser 2 4 0.00000000033832
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206060_1.5nF
*******
.subckt 0603_885012206061_2.2nF 1 2
Rser 1 3 0.12731
Lser 2 4 0.00000000032293
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012206061_2.2nF
*******
.subckt 0603_885012206062_3.3nF 1 2
Rser 1 3 0.09865
Lser 2 4 0.0000000003316
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206062_3.3nF
*******
.subckt 0603_885012206063_4.7nF 1 2
Rser 1 3 0.08147
Lser 2 4 0.0000000002893
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206063_4.7nF
*******
.subckt 0603_885012206064_6.8nF 1 2
Rser 1 3 0.08487
Lser 2 4 0.00000000036849
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206064_6.8nF
*******
.subckt 0603_885012206065_10nF 1 2
Rser 1 3 0.05893
Lser 2 4 0.00000000037916
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206065_10nF
*******
.subckt 0603_885012206066_15nF 1 2
Rser 1 3 0.0473
Lser 2 4 0.00000000030093
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0603_885012206066_15nF
*******
.subckt 0603_885012206067_22nF 1 2
Rser 1 3 0.03101
Lser 2 4 0.00000000028048
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885012206067_22nF
*******
.subckt 0603_885012206068_33nF 1 2
Rser 1 3 0.0232
Lser 2 4 0.00000000033089
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0603_885012206068_33nF
*******
.subckt 0603_885012206069_47nF 1 2
Rser 1 3 0.01832
Lser 2 4 0.0000000002418
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0603_885012206069_47nF
*******
.subckt 0603_885012206070_68nF 1 2
Rser 1 3 0.01712
Lser 2 4 0.00000000030682
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0603_885012206070_68nF
*******
.subckt 0603_885012206071_100nF 1 2
Rser 1 3 0.025
Lser 2 4 0.0000000008
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206071_100nF
*******
.subckt 0603_885012206072_150nF 1 2
Rser 1 3 0.0149181934238
Lser 2 4 3.31198563E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0603_885012206072_150nF
*******
.subckt 0603_885012206073_220nF 1 2
Rser 1 3 0.0109800094243
Lser 2 4 4.08100466E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012206073_220nF
*******
.subckt 0603_885012206074_330nF 1 2
Rser 1 3 0.0118150527569
Lser 2 4 4.48623546E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012206074_330nF
*******
.subckt 0603_885012206075_470nF 1 2
Rser 1 3 0.0100816359349
Lser 2 4 4.14055319E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012206075_470nF
*******
.subckt 0603_885012206076_1uF 1 2
Rser 1 3 0.0073448307676
Lser 2 4 4.75503387E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0603_885012206076_1uF
*******
.subckt 0603_885012206071R_100nF 1 2
Rser 1 3 0.0189365521551
Lser 2 4 4.42668552E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206071R_100nF
*******
.subckt 0603_885012206075R_470nF 1 2
Rser 1 3 0.0100816359349
Lser 2 4 4.14055319E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0603_885012206075R_470nF
*******
.subckt 0805_885012007026_3.3pF 1 2
Rser 1 3 0.407676004204
Lser 2 4 4.49191488E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0805_885012007026_3.3pF
*******
.subckt 0805_885012007027_6.8pF 1 2
Rser 1 3 0.359480200218
Lser 2 4 4.5722648E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0805_885012007027_6.8pF
*******
.subckt 0805_885012007028_10pF 1 2
Rser 1 3 0.366485482781
Lser 2 4 5.23706793E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0805_885012007028_10pF
*******
.subckt 0805_885012007029_15pF 1 2
Rser 1 3 0.322140605571
Lser 2 4 5.33099942E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007029_15pF
*******
.subckt 0805_885012007030_22pF 1 2
Rser 1 3 0.337501541959
Lser 2 4 6.08362599E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0805_885012007030_22pF
*******
.subckt 0805_885012007031_33pF 1 2
Rser 1 3 0.266905660637
Lser 2 4 5.7081292E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007031_33pF
*******
.subckt 0805_885012007032_47pF 1 2
Rser 1 3 0.224971777912
Lser 2 4 5.50463607E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885012007032_47pF
*******
.subckt 0805_885012007033_68pF 1 2
Rser 1 3 0.188385732986
Lser 2 4 4.4496757E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0805_885012007033_68pF
*******
.subckt 0805_885012007034_100pF 1 2
Rser 1 3 0.118679326168
Lser 2 4 2.41991847E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007034_100pF
*******
.subckt 0805_885012007035_150pF 1 2
Rser 1 3 0.135556605699
Lser 2 4 4.3127146E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007035_150pF
*******
.subckt 0805_885012007036_220pF 1 2
Rser 1 3 0.115723179071
Lser 2 4 4.36175568E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012007036_220pF
*******
.subckt 0805_885012007037_330pF 1 2
Rser 1 3 0.0911424032195
Lser 2 4 4.34684674E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007037_330pF
*******
.subckt 0805_885012007038_470pF 1 2
Rser 1 3 0.0888157768288
Lser 2 4 4.59255914E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007038_470pF
*******
.subckt 0805_885012007039_680pF 1 2
Rser 1 3 0.0750121415022
Lser 2 4 4.46094349E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012007039_680pF
*******
.subckt 0805_885012007040_1nF 1 2
Rser 1 3 0.0506576337129
Lser 2 4 2.60606775E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007040_1nF
*******
.subckt 0805_885012007041_1.5nF 1 2
Rser 1 3 0.0403337213614
Lser 2 4 2.897145E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012007041_1.5nF
*******
.subckt 0805_885012007042_2.2nF 1 2
Rser 1 3 0.0313104040283
Lser 2 4 2.67647833E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012007042_2.2nF
*******
.subckt 0805_885012007043_3.3nF 1 2
Rser 1 3 0.0278586078187
Lser 2 4 3.06758727E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012007043_3.3nF
*******
.subckt 0805_885012007044_4.7nF 1 2
Rser 1 3 0.0125481242528
Lser 2 4 1.0825546E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012007044_4.7nF
*******
.subckt 0805_885012107015_1uF 1 2
Rser 1 3 0.00799934804354
Lser 2 4 2.55135429E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885012107015_1uF
*******
.subckt 0805_885012107016_2.2uF 1 2
Rser 1 3 0.00497944150425
Lser 2 4 2.69972955E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012107016_2.2uF
*******
.subckt 0805_885012107017_3.3uF 1 2
Rser 1 3 0.0041415980008
Lser 2 4 2.72087954E-10
C1 3 4 0.0000033
Rpar 3 4 30000000
.ends 0805_885012107017_3.3uF
*******
.subckt 0805_885012107018_4.7uF 1 2
Rser 1 3 0.00349429730952
Lser 2 4 2.52123218E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 0805_885012107018_4.7uF
*******
.subckt 0805_885012207054_100pF 1 2
Rser 1 3 0.90625
Lser 2 4 0.00000000029357
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207054_100pF
*******
.subckt 0805_885012207055_150pF 1 2
Rser 1 3 0.70433
Lser 2 4 0.00000000030352
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012207055_150pF
*******
.subckt 0805_885012207056_220pF 1 2
Rser 1 3 0.48805
Lser 2 4 0.00000000027764
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012207056_220pF
*******
.subckt 0805_885012207057_330pF 1 2
Rser 1 3 0.44753
Lser 2 4 0.00000000032997
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012207057_330pF
*******
.subckt 0805_885012207058_470pF 1 2
Rser 1 3 0.32032
Lser 2 4 0.0000000002982
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207058_470pF
*******
.subckt 0805_885012207059_680pF 1 2
Rser 1 3 0.25951
Lser 2 4 0.00000000036777
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012207059_680pF
*******
.subckt 0805_885012207060_1nF 1 2
Rser 1 3 0.20128
Lser 2 4 0.00000000029022
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207060_1nF
*******
.subckt 0805_885012207061_1.5nF 1 2
Rser 1 3 0.15833
Lser 2 4 0.00000000037277
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207061_1.5nF
*******
.subckt 0805_885012207062_2.2nF 1 2
Rser 1 3 0.11878
Lser 2 4 0.00000000036877
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012207062_2.2nF
*******
.subckt 0805_885012207063_3.3nF 1 2
Rser 1 3 0.10404
Lser 2 4 0.00000000034071
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207063_3.3nF
*******
.subckt 0805_885012207064_4.7nF 1 2
Rser 1 3 0.07475
Lser 2 4 0.00000000024317
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012207064_4.7nF
*******
.subckt 0805_885012207065_6.8nF 1 2
Rser 1 3 0.08276
Lser 2 4 0.00000000032015
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0805_885012207065_6.8nF
*******
.subckt 0805_885012207066_10nF 1 2
Rser 1 3 0.06408
Lser 2 4 0.0000000002943
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207066_10nF
*******
.subckt 0805_885012207067_15nF 1 2
Rser 1 3 0.05208
Lser 2 4 0.00000000031399
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0805_885012207067_15nF
*******
.subckt 0805_885012207068_22nF 1 2
Rser 1 3 0.0486328028818
Lser 2 4 0.00000000041
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0805_885012207068_22nF
*******
.subckt 0805_885012207069_33nF 1 2
Rser 1 3 0.0330484373884
Lser 2 4 0.00000000041
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0805_885012207069_33nF
*******
.subckt 0805_885012207070_47nF 1 2
Rser 1 3 0.0298909488495
Lser 2 4 0.00000000038
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0805_885012207070_47nF
*******
.subckt 0805_885012207071_68nF 1 2
Rser 1 3 0.0247
Lser 2 4 0.00000000027034
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0805_885012207071_68nF
*******
.subckt 0805_885012207072_100nF 1 2
Rser 1 3 0.0172819633028
Lser 2 4 0.00000000035
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207072_100nF
*******
.subckt 0805_885012207073_150nF 1 2
Rser 1 3 0.0145783171748
Lser 2 4 0.00000000035
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0805_885012207073_150nF
*******
.subckt 0805_885012207074_220nF 1 2
Rser 1 3 0.0111697818844
Lser 2 4 0.00000000042
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885012207074_220nF
*******
.subckt 0805_885012207075_330nF 1 2
Rser 1 3 0.00939488017121
Lser 2 4 0.000000000283
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885012207075_330nF
*******
.subckt 0805_885012207076_470nF 1 2
Rser 1 3 0.00781019032257
Lser 2 4 0.00000000049
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0805_885012207076_470nF
*******
.subckt 0805_885012207077_680nF 1 2
Rser 1 3 0.00783503615977
Lser 2 4 0.00000000053
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 0805_885012207077_680nF
*******
.subckt 0805_885012207078_1uF 1 2
Rser 1 3 0.00804838198988
Lser 2 4 2.69843792E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0805_885012207078_1uF
*******
.subckt 0805_885012207079_2.2uF 1 2
Rser 1 3 0.00468718250549
Lser 2 4 2.80891331E-10
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 0805_885012207079_2.2uF
*******
.subckt 0805_885012107019_22uF 1 2
Rser 1 3 0.006
Lser 2 4 0.000000000834
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 0805_885012107019_22uF
*******
.subckt 0805_885012107027_10uF 1 2
Rser 1 3 0.007
Lser 2 4 0.0000000009
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 0805_885012107027_10uF
*******
.subckt 1206_885012008019_10pF 1 2
Rser 1 3 0.391301643484
Lser 2 4 5.83813577E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1206_885012008019_10pF
*******
.subckt 1206_885012008020_33pF 1 2
Rser 1 3 0.254333105283
Lser 2 4 4.78321618E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 1206_885012008020_33pF
*******
.subckt 1206_885012008021_47pF 1 2
Rser 1 3 0.233708673806
Lser 2 4 4.88472845E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885012008021_47pF
*******
.subckt 1206_885012008022_68pF 1 2
Rser 1 3 0.199591933016
Lser 2 4 4.68378192E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 1206_885012008022_68pF
*******
.subckt 1206_885012008023_100pF 1 2
Rser 1 3 0.15525411437
Lser 2 4 4.47352225E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008023_100pF
*******
.subckt 1206_885012008024_330pF 1 2
Rser 1 3 0.0916318679708
Lser 2 4 3.11969377E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012008024_330pF
*******
.subckt 1206_885012008025_470pF 1 2
Rser 1 3 0.106551883888
Lser 2 4 4.30008474E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012008025_470pF
*******
.subckt 1206_885012008026_1nF 1 2
Rser 1 3 0.0693861515837
Lser 2 4 4.13253027E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012008026_1nF
*******
.subckt 1206_885012008027_2.2nF 1 2
Rser 1 3 0.0393800076857
Lser 2 4 5.03985839E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012008027_2.2nF
*******
.subckt 1206_885012008028_4.7nF 1 2
Rser 1 3 0.0260664466932
Lser 2 4 4.4983761E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012008028_4.7nF
*******
.subckt 1206_885012008029_6.8nF 1 2
Rser 1 3 0.0469294057584
Lser 2 4 4.43201944E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008029_6.8nF
*******
.subckt 1206_885012008030_10nF 1 2
Rser 1 3 0.0261734331747
Lser 2 4 5.33952576E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008030_10nF
*******
.subckt 1206_885012108019_2.2uF 1 2
Rser 1 3 0.00474329771021
Lser 2 4 5.16937352E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012108019_2.2uF
*******
.subckt 1206_885012108020_4.7uF 1 2
Rser 1 3 0.00541345635951
Lser 2 4 5.0768239E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1206_885012108020_4.7uF
*******
.subckt 1206_885012108021_10uF 1 2
Rser 1 3 0.00349318752029
Lser 2 4 6.43774867E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012108021_10uF
*******
.subckt 1206_885012208042_220pF 1 2
Rser 1 3 0.58352
Lser 2 4 0.00000000032083
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012208042_220pF
*******
.subckt 1206_885012208043_330pF 1 2
Rser 1 3 0.50009
Lser 2 4 0.00000000035086
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012208043_330pF
*******
.subckt 1206_885012208044_470pF 1 2
Rser 1 3 0.35551
Lser 2 4 0.0000000004724
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208044_470pF
*******
.subckt 1206_885012208045_680pF 1 2
Rser 1 3 0.32598
Lser 2 4 0.0000000006527
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012208045_680pF
*******
.subckt 1206_885012208046_1nF 1 2
Rser 1 3 0.23112
Lser 2 4 0.00000000050124
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208046_1nF
*******
.subckt 1206_885012208047_1.5nF 1 2
Rser 1 3 0.17032
Lser 2 4 0.00000000040983
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012208047_1.5nF
*******
.subckt 1206_885012208048_2.2nF 1 2
Rser 1 3 0.11761
Lser 2 4 0.00000000058541
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012208048_2.2nF
*******
.subckt 1206_885012208049_3.3nF 1 2
Rser 1 3 0.12683
Lser 2 4 0.00000000044431
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012208049_3.3nF
*******
.subckt 1206_885012208050_4.7nF 1 2
Rser 1 3 0.07742
Lser 2 4 0.00000000042481
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208050_4.7nF
*******
.subckt 1206_885012208051_6.8nF 1 2
Rser 1 3 0.0893088703811
Lser 2 4 5.44959228E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012208051_6.8nF
*******
.subckt 1206_885012208052_10nF 1 2
Rser 1 3 0.355515780687
Lser 2 4 4.90239917E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208052_10nF
*******
.subckt 1206_885012208053_15nF 1 2
Rser 1 3 0.05086
Lser 2 4 0.00000000064474
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1206_885012208053_15nF
*******
.subckt 1206_885012208054_22nF 1 2
Rser 1 3 0.04388
Lser 2 4 0.00000000043595
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1206_885012208054_22nF
*******
.subckt 1206_885012208055_33nF 1 2
Rser 1 3 0.05974
Lser 2 4 0.00000000046935
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1206_885012208055_33nF
*******
.subckt 1206_885012208056_47nF 1 2
Rser 1 3 0.05553
Lser 2 4 0.00000000049393
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1206_885012208056_47nF
*******
.subckt 1206_885012208057_68nF 1 2
Rser 1 3 0.03879
Lser 2 4 0.00000000044546
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 1206_885012208057_68nF
*******
.subckt 1206_885012208058_100nF 1 2
Rser 1 3 0.0232208356231
Lser 2 4 5.59299026E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885012208058_100nF
*******
.subckt 1206_885012208059_150nF 1 2
Rser 1 3 0.0179362383614
Lser 2 4 5.89126458E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1206_885012208059_150nF
*******
.subckt 1206_885012208060_220nF 1 2
Rser 1 3 0.0124482582844
Lser 2 4 5.568771E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1206_885012208060_220nF
*******
.subckt 1206_885012208061_330nF 1 2
Rser 1 3 0.0123070322618
Lser 2 4 7.16267872E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1206_885012208061_330nF
*******
.subckt 1206_885012208062_470nF 1 2
Rser 1 3 0.0100846165597
Lser 2 4 7.45549291E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1206_885012208062_470nF
*******
.subckt 1206_885012208063_680nF 1 2
Rser 1 3 0.00806863562842
Lser 2 4 7.09595993E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1206_885012208063_680nF
*******
.subckt 1206_885012208064_1uF 1 2
Rser 1 3 0.00633398843665
Lser 2 4 7.50258152E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885012208064_1uF
*******
.subckt 1206_885012208065_1.5uF 1 2
Rser 1 3 0.00655648262409
Lser 2 4 8.57454998E-10
C1 3 4 0.0000015
Rpar 3 4 300000000
.ends 1206_885012208065_1.5uF
*******
.subckt 1206_885012208066_2.2uF 1 2
Rser 1 3 0.00520440828302
Lser 2 4 7.87876644E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1206_885012208066_2.2uF
*******
.subckt 1206_885012208067_3.3uF 1 2
Rser 1 3 0.00537091922132
Lser 2 4 8.20379233E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1206_885012208067_3.3uF
*******
.subckt 1206_885012208068_4.7uF 1 2
Rser 1 3 0.00336451412099
Lser 2 4 7.97503693E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1206_885012208068_4.7uF
*******
.subckt 1206_885012208069_10uF 1 2
Rser 1 3 0.0039007012861
Lser 2 4 0.00000000055
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012208069_10uF
*******
.subckt 1210_885012009002_1nF 1 2
Rser 1 3 0.0526199422099
Lser 2 4 2.28139939E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885012009002_1nF
*******
.subckt 1210_885012009003_2.2nF 1 2
Rser 1 3 0.236239384732
Lser 2 4 2.48857755E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1210_885012009003_2.2nF
*******
.subckt 1210_885012009004_4.7nF 1 2
Rser 1 3 0.0889145917519
Lser 2 4 2.66275966E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1210_885012009004_4.7nF
*******
.subckt 1210_885012009005_6.8nF 1 2
Rser 1 3 0.0165690812867
Lser 2 4 2.56210234E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1210_885012009005_6.8nF
*******
.subckt 1210_885012009006_15nF 1 2
Rser 1 3 0.0164446208365
Lser 2 4 3.024777E-10
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1210_885012009006_15nF
*******
.subckt 1210_885012109012_4.7uF 1 2
Rser 1 3 0.0033906445918
Lser 2 4 3.01326093E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012109012_4.7uF
*******
.subckt 1210_885012109013_10uF 1 2
Rser 1 3 0.00241697975791
Lser 2 4 8.77086276E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1210_885012109013_10uF
*******
.subckt 1210_885012109014_22uF 1 2
Rser 1 3 0.00268514753558
Lser 2 4 9.0689132E-10
C1 3 4 0.000022
Rpar 3 4 2000000
.ends 1210_885012109014_22uF
*******
.subckt 1210_885012109015_22uF 1 2
Rser 1 3 0.00734474129923
Lser 2 4 1.236549611E-09
C1 3 4 0.000022
Rpar 3 4 5000000
.ends 1210_885012109015_22uF
*******
.subckt 1210_885012209015_1nF 1 2
Rser 1 3 0.23064
Lser 2 4 0.00000000009004
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885012209015_1nF
*******
.subckt 1210_885012209016_2.2nF 1 2
Rser 1 3 0.15
Lser 2 4 0.0000000009
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1210_885012209016_2.2nF
*******
.subckt 1210_885012209017_10nF 1 2
Rser 1 3 0.07411
Lser 2 4 0.00000000018051
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1210_885012209017_10nF
*******
.subckt 1210_885012209018_22nF 1 2
Rser 1 3 0.06131
Lser 2 4 0.00000000020837
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1210_885012209018_22nF
*******
.subckt 1210_885012209019_100nF 1 2
Rser 1 3 0.0209574310072
Lser 2 4 5.49171232E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1210_885012209019_100nF
*******
.subckt 1210_885012209020_220nF 1 2
Rser 1 3 0.0109918196754
Lser 2 4 5.14177759E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1210_885012209020_220nF
*******
.subckt 1210_885012209021_330nF 1 2
Rser 1 3 0.00972375707294
Lser 2 4 5.4771949E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1210_885012209021_330nF
*******
.subckt 1210_885012209022_470nF 1 2
Rser 1 3 0.00740093895541
Lser 2 4 5.16300103E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1210_885012209022_470nF
*******
.subckt 1210_885012209023_680nF 1 2
Rser 1 3 0.00560873026626
Lser 2 4 5.62947674E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1210_885012209023_680nF
*******
.subckt 1210_885012209024_1uF 1 2
Rser 1 3 0.00434521559376
Lser 2 4 3.4952573E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209024_1uF
*******
.subckt 1210_885012209025_2.2uF 1 2
Rser 1 3 0.003755566195
Lser 2 4 4.76192409E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1210_885012209025_2.2uF
*******
.subckt 1210_885012209026_3.3uF 1 2
Rser 1 3 0.0037725139254
Lser 2 4 4.43584901E-10
C1 3 4 0.0000033
Rpar 3 4 200000000
.ends 1210_885012209026_3.3uF
*******
.subckt 1210_885012209027_4.7uF 1 2
Rser 1 3 0.00334303070776
Lser 2 4 4.2432524E-10
C1 3 4 0.0000047
Rpar 3 4 100000000
.ends 1210_885012209027_4.7uF
*******
.subckt 1210_885012209028_10uF 1 2
Rser 1 3 0.0026086390311
Lser 2 4 8.94000611E-10
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 1210_885012209028_10uF
*******
.subckt 1210_885012209074_22uF 1 2
Rser 1 3 0.0043
Lser 2 4 0.000000001
C1 3 4 0.000022
Rpar 3 4 5000000
.ends 1210_885012209074_22uF
*******
.subckt 1812_885012010003_10nF 1 2
Rser 1 3 0.035610362113
Lser 2 4 2.40113972E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012010003_10nF
*******
.subckt 1812_885012010004_33nF 1 2
Rser 1 3 0.0120609525555
Lser 2 4 3.8469537E-10
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1812_885012010004_33nF
*******
.subckt 1812_885012210005_4.7nF 1 2
Rser 1 3 0.0828
Lser 2 4 0.00000000018862
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1812_885012210005_4.7nF
*******
.subckt 1812_885012210006_10nF 1 2
Rser 1 3 0.07693
Lser 2 4 0.00000000053548
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012210006_10nF
*******
.subckt 1812_885012210007_47nF 1 2
Rser 1 3 0.03468
Lser 2 4 0.00000000076842
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1812_885012210007_47nF
*******
.subckt 1812_885012210008_100nF 1 2
Rser 1 3 0.037008688888
Lser 2 4 6.73793576E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1812_885012210008_100nF
*******
.subckt 1812_885012210009_330nF 1 2
Rser 1 3 0.01427157177
Lser 2 4 4.80558989E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1812_885012210009_330nF
*******
.subckt 1812_885012210010_470nF 1 2
Rser 1 3 0.00985565119595
Lser 2 4 4.00753105E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1812_885012210010_470nF
*******
.subckt 1812_885012210011_680nF 1 2
Rser 1 3 0.00784524987635
Lser 2 4 4.30816782E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1812_885012210011_680nF
*******
.subckt 1812_885012210012_1uF 1 2
Rser 1 3 0.014
Lser 2 4 0.000000001
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1812_885012210012_1uF
*******
.subckt 2220_885012214004_10uF 1 2
Rser 1 3 0.003
Lser 2 4 0.0000000012
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 2220_885012214004_10uF
*******
