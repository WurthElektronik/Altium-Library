**************************************************
* Manufacturer:          Würth Elektronik 
* Kinds:                 SMT Power Inductor
* Matchcode:             WE-LHMI
* Library Type:          LTspice
* Version:               rev23a
* Created/modified by:   Ella
* Date and Time:         8/14/2023
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2023 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 1040_74437368010_1u  1 2
Rp 1 2 941.74
Cp 1 2 13.7p
Rs 1 N3 0.003
L1 N3 2 0.91u
.ends 1040_74437368010_1u 
*******
.subckt 1040_74437368022_2.2u  1 2
Rp 1 2 1611.67
Cp 1 2 18.93p
Rs 1 N3 0.0065
L1 N3 2 1.82u
.ends 1040_74437368022_2.2u 
*******
.subckt 1040_74437368033_3.3u  1 2
Rp 1 2 2310.37
Cp 1 2 18.43p
Rs 1 N3 0.0108
L1 N3 2 2.84u
.ends 1040_74437368033_3.3u 
*******
.subckt 1040_74437368039_3.9u  1 2
Rp 1 2 5533
Cp 1 2 24.83p
Rs 1 N3 0.0126
L1 N3 2 3.9u
.ends 1040_74437368039_3.9u 
*******
.subckt 1040_74437368047_4.7u  1 2
Rp 1 2 2644.46
Cp 1 2 22.64p
Rs 1 N3 0.015
L1 N3 2 3.98u
.ends 1040_74437368047_4.7u 
*******
.subckt 1040_74437368056_5.6u  1 2
Rp 1 2 2629
Cp 1 2 25.756p
Rs 1 N3 0.0176
L1 N3 2 5.6u
.ends 1040_74437368056_5.6u 
*******
.subckt 1040_74437368068_6.8u  1 2
Rp 1 2 3702.85
Cp 1 2 24.69p
Rs 1 N3 0.0175
L1 N3 2 6.38u
.ends 1040_74437368068_6.8u 
*******
.subckt 1040_74437368100_10u  1 2
Rp 1 2 5143.82666666667
Cp 1 2 18.6066666666667p
Rs 1 N3 0.027
L1 N3 2 8.6u
.ends 1040_74437368100_10u 
*******
.subckt 1040_74437368150_15u  1 2
Rp 1 2 10500
Cp 1 2 26.338p
Rs 1 N3 0.04
L1 N3 2 14.48u
.ends 1040_74437368150_15u 
*******
.subckt 1040_74437368220_22u  1 2
Rp 1 2 18986
Cp 1 2 23.505p
Rs 1 N3 0.064
L1 N3 2 18.99u
.ends 1040_74437368220_22u 
*******
.subckt 1040_74437368330_33u  1 2
Rp 1 2 30592
Cp 1 2 25.532p
Rs 1 N3 0.092
L1 N3 2 30.95u
.ends 1040_74437368330_33u 
*******
.subckt 1040_74437368470_47u  1 2
Rp 1 2 20405
Cp 1 2 22.1p
Rs 1 N3 0.145
L1 N3 2 47u
.ends 1040_74437368470_47u 
*******
.subckt 1040_744373680022_0.22u  1 2
Rp 1 2 327.73
Cp 1 2 5.25p
Rs 1 N3 0.0008
L1 N3 2 0.2u
.ends 1040_744373680022_0.22u 
*******
.subckt 1040_744373680036_0.36u  1 2
Rp 1 2 376.64
Cp 1 2 8.58p
Rs 1 N3 0.00105
L1 N3 2 0.29u
.ends 1040_744373680036_0.36u 
*******
.subckt 1040_744373680039_0.39u  1 2
Rp 1 2 392.21
Cp 1 2 7.35p
Rs 1 N3 0.0011
L1 N3 2 0.32u
.ends 1040_744373680039_0.39u 
*******
.subckt 1040_744373680045_0.45u  1 2
Rp 1 2 555.32
Cp 1 2 8.87p
Rs 1 N3 0.0013
L1 N3 2 0.45u
.ends 1040_744373680045_0.45u 
*******
.subckt 1040_744373680056_0.56u  1 2
Rp 1 2 509.43
Cp 1 2 10.4p
Rs 1 N3 0.0016
L1 N3 2 0.5u
.ends 1040_744373680056_0.56u 
*******
.subckt 1040_744373680068_0.68u  1 2
Rp 1 2 509.43
Cp 1 2 10.4p
Rs 1 N3 0.0024
L1 N3 2 0.68u
.ends 1040_744373680068_0.68u 
*******
.subckt 1335_74437377010_1u  1 2
Rp 1 2 731.66
Cp 1 2 15.61p
Rs 1 N3 0.0027
L1 N3 2 0.97u
.ends 1335_74437377010_1u 
*******
.subckt 1335_74437377015_1.5u  1 2
Rp 1 2 1636.07
Cp 1 2 21.23p
Rs 1 N3 0.0047
L1 N3 2 1.39u
.ends 1335_74437377015_1.5u 
*******
.subckt 1335_74437377022_2.2u  1 2
Rp 1 2 2241
Cp 1 2 23.99p
Rs 1 N3 0.0072
L1 N3 2 2.18u
.ends 1335_74437377022_2.2u 
*******
.subckt 1335_74437377033_3.3u  1 2
Rp 1 2 2736.47
Cp 1 2 30.65p
Rs 1 N3 0.009
L1 N3 2 2.89u
.ends 1335_74437377033_3.3u 
*******
.subckt 1335_74437377047_4.7u  1 2
Rp 1 2 2277.33
Cp 1 2 34.92p
Rs 1 N3 0.013
L1 N3 2 4.3u
.ends 1335_74437377047_4.7u 
*******
.subckt 1335_744373770022_0.22u  1 2
Rp 1 2 270.32
Cp 1 2 7.64p
Rs 1 N3 0.00075
L1 N3 2 0.21u
.ends 1335_744373770022_0.22u 
*******
.subckt 1335_744373770033_0.33u  1 2
Rp 1 2 321.42
Cp 1 2 8.3p
Rs 1 N3 0.00088
L1 N3 2 0.31u
.ends 1335_744373770033_0.33u 
*******
.subckt 1335_744373770047_0.47u  1 2
Rp 1 2 542.84
Cp 1 2 9.8p
Rs 1 N3 0.00132
L1 N3 2 0.46u
.ends 1335_744373770047_0.47u 
*******
.subckt 1335_744373770056_0.56u  1 2
Rp 1 2 581.77
Cp 1 2 13.88p
Rs 1 N3 0.0014
L1 N3 2 0.54u
.ends 1335_744373770056_0.56u 
*******
.subckt 1335_744373770068_0.68u  1 2
Rp 1 2 817.29
Cp 1 2 15.04p
Rs 1 N3 0.0018
L1 N3 2 0.66u
.ends 1335_744373770068_0.68u 
*******
.subckt 1365_744373965010_1u  1 2
Rp 1 2 1359
Cp 1 2 15.41p
Rs 1 N3 0.0019
L1 N3 2 1u
.ends 1365_744373965010_1u 
*******
.subckt 1365_744373965015_1.5u  1 2
Rp 1 2 1358
Cp 1 2 19.52p
Rs 1 N3 0.0023
L1 N3 2 1.5u
.ends 1365_744373965015_1.5u 
*******
.subckt 1365_744373965022_2.2u  1 2
Rp 1 2 1941
Cp 1 2 25.74p
Rs 1 N3 0.0032
L1 N3 2 2.2u
.ends 1365_744373965022_2.2u 
*******
.subckt 1365_744373965033_3.3u  1 2
Rp 1 2 6035
Cp 1 2 20.92p
Rs 1 N3 0.0057
L1 N3 2 3.3u
.ends 1365_744373965033_3.3u 
*******
.subckt 1365_744373965047_4.7u  1 2
Rp 1 2 6592
Cp 1 2 27.48p
Rs 1 N3 0.0065
L1 N3 2 4.7u
.ends 1365_744373965047_4.7u 
*******
.subckt 1365_744373965056_5.6u  1 2
Rp 1 2 6916
Cp 1 2 27.15p
Rs 1 N3 0.0083
L1 N3 2 5.6u
.ends 1365_744373965056_5.6u 
*******
.subckt 1365_744373965068_6.8u  1 2
Rp 1 2 8283
Cp 1 2 29.96p
Rs 1 N3 0.0092
L1 N3 2 6.8u
.ends 1365_744373965068_6.8u 
*******
.subckt 1365_744373965100_10u  1 2
Rp 1 2 4157
Cp 1 2 40.93p
Rs 1 N3 0.0106
L1 N3 2 10u
.ends 1365_744373965100_10u 
*******
.subckt 1365_744373965101_100u  1 2
Rp 1 2 12541
Cp 1 2 44.96p
Rs 1 N3 0.1408
L1 N3 2 100u
.ends 1365_744373965101_100u 
*******
.subckt 1365_744373965120_12u  1 2
Rp 1 2 5228
Cp 1 2 39.71p
Rs 1 N3 0.0178
L1 N3 2 12u
.ends 1365_744373965120_12u 
*******
.subckt 1365_744373965150_15u  1 2
Rp 1 2 6124
Cp 1 2 29.55p
Rs 1 N3 0.0244
L1 N3 2 15u
.ends 1365_744373965150_15u 
*******
.subckt 1365_744373965220_22u  1 2
Rp 1 2 7428
Cp 1 2 37p
Rs 1 N3 0.0345
L1 N3 2 22u
.ends 1365_744373965220_22u 
*******
.subckt 1365_744373965330_33u  1 2
Rp 1 2 9823
Cp 1 2 39.64p
Rs 1 N3 0.0487
L1 N3 2 33u
.ends 1365_744373965330_33u 
*******
.subckt 1365_744373965470_47u  1 2
Rp 1 2 8647
Cp 1 2 40.74p
Rs 1 N3 0.0746
L1 N3 2 47u
.ends 1365_744373965470_47u 
*******
.subckt 1365_7443739650022_0.22u  1 2
Rp 1 2 439.566
Cp 1 2 10.36p
Rs 1 N3 0.00051
L1 N3 2 0.22u
.ends 1365_7443739650022_0.22u 
*******
.subckt 1365_7443739650033_0.33u  1 2
Rp 1 2 531.88
Cp 1 2 14.12p
Rs 1 N3 0.00064
L1 N3 2 0.33u
.ends 1365_7443739650033_0.33u 
*******
.subckt 1365_7443739650047_0.47u  1 2
Rp 1 2 698.73
Cp 1 2 15.7p
Rs 1 N3 0.00092
L1 N3 2 0.47u
.ends 1365_7443739650047_0.47u 
*******
.subckt 1365_7443739650056_0.56u  1 2
Rp 1 2 357.47
Cp 1 2 17.34p
Rs 1 N3 0.00111
L1 N3 2 0.56u
.ends 1365_7443739650056_0.56u 
*******
.subckt 1365_7443739650068_0.68u  1 2
Rp 1 2 384.64
Cp 1 2 15.95p
Rs 1 N3 0.0012
L1 N3 2 0.68u
.ends 1365_7443739650068_0.68u 
*******
.subckt 4012_74437321010_1u  1 2
Rp 1 2 2449.262983768
Cp 1 2 3.62591534p
Rs 1 N3 0.041
L1 N3 2 0.85u
.ends 4012_74437321010_1u 
*******
.subckt 4012_74437321015_1.5u  1 2
Rp 1 2 3509.095675436
Cp 1 2 4.622831186p
Rs 1 N3 0.055
L1 N3 2 1.46u
.ends 4012_74437321015_1.5u 
*******
.subckt 4012_74437321022_2.2u  1 2
Rp 1 2 5186.32963784
Cp 1 2 3.9005875664p
Rs 1 N3 0.0692
L1 N3 2 1.98u
.ends 4012_74437321022_2.2u 
*******
.subckt 4012_74437321033_3.3u  1 2
Rp 1 2 6592.331864912
Cp 1 2 5.2925305872p
Rs 1 N3 0.084
L1 N3 2 3.09u
.ends 4012_74437321033_3.3u 
*******
.subckt 4012_74437321047_4.7u  1 2
Rp 1 2 8647.359812636
Cp 1 2 5.2991188784p
Rs 1 N3 0.128
L1 N3 2 4.44u
.ends 4012_74437321047_4.7u 
*******
.subckt 4012_74437321056_5.6u  1 2
Rp 1 2 9952.654835202
Cp 1 2 5.7131337644p
Rs 1 N3 0.18
L1 N3 2 5.64u
.ends 4012_74437321056_5.6u 
*******
.subckt 4012_74437321068_6.8u  1 2
Rp 1 2 11916.18781332
Cp 1 2 5.7684705248p
Rs 1 N3 0.3
L1 N3 2 7u
.ends 4012_74437321068_6.8u 
*******
.subckt 4012_74437321082_8.2u  1 2
Rp 1 2 14407.6610493
Cp 1 2 5.3210721894p
Rs 1 N3 0.313
L1 N3 2 8.17u
.ends 4012_74437321082_8.2u 
*******
.subckt 4012_74437321100_10u  1 2
Rp 1 2 17155.04252754
Cp 1 2 5.3301573364p
Rs 1 N3 0.41
L1 N3 2 9.27u
.ends 4012_74437321100_10u 
*******
.subckt 4012_744373210010_0.1u  1 2
Rp 1 2 361.4225009824
Cp 1 2 2.3572271464p
Rs 1 N3 0.0043
L1 N3 2 0.082u
.ends 4012_744373210010_0.1u 
*******
.subckt 4012_744373210022_0.22u  1 2
Rp 1 2 620.2025012388
Cp 1 2 2.9064357274p
Rs 1 N3 0.0066
L1 N3 2 0.17u
.ends 4012_744373210022_0.22u 
*******
.subckt 4012_744373210047_0.47u  1 2
Rp 1 2 1209.327994442
Cp 1 2 3.698166362p
Rs 1 N3 0.018
L1 N3 2 0.45u
.ends 4012_744373210047_0.47u 
*******
.subckt 4020_74437324010_1u  1 2
Rp 1 2 1017.16
Cp 1 2 4.16p
Rs 1 N3 0.022
L1 N3 2 0.79u
.ends 4020_74437324010_1u 
*******
.subckt 4020_74437324012_1.2u  1 2
Rp 1 2 1114.36
Cp 1 2 5.1p
Rs 1 N3 0.025
L1 N3 2 1.02u
.ends 4020_74437324012_1.2u 
*******
.subckt 4020_74437324015_1.5u  1 2
Rp 1 2 1434.01
Cp 1 2 4.71p
Rs 1 N3 0.0348
L1 N3 2 1.33u
.ends 4020_74437324015_1.5u 
*******
.subckt 4020_74437324022_2.2u  1 2
Rp 1 2 2011.68
Cp 1 2 5.56p
Rs 1 N3 0.051
L1 N3 2 1.92u
.ends 4020_74437324022_2.2u 
*******
.subckt 4020_74437324033_3.3u  1 2
Rp 1 2 2663.25
Cp 1 2 5.59p
Rs 1 N3 0.069
L1 N3 2 2.98u
.ends 4020_74437324033_3.3u 
*******
.subckt 4020_74437324047_4.7u  1 2
Rp 1 2 3800.41
Cp 1 2 6.26p
Rs 1 N3 0.095
L1 N3 2 4.42u
.ends 4020_74437324047_4.7u 
*******
.subckt 4020_74437324056_5.6u  1 2
Rp 1 2 4331.66
Cp 1 2 6.06p
Rs 1 N3 0.12
L1 N3 2 4.94u
.ends 4020_74437324056_5.6u 
*******
.subckt 4020_74437324068_6.8u  1 2
Rp 1 2 4993.38
Cp 1 2 5.8p
Rs 1 N3 0.15
L1 N3 2 5.31u
.ends 4020_74437324068_6.8u 
*******
.subckt 4020_74437324082_8.2u  1 2
Rp 1 2 4933.23
Cp 1 2 6.207p
Rs 1 N3 0.158
L1 N3 2 7.91u
.ends 4020_74437324082_8.2u 
*******
.subckt 4020_74437324100_10u  1 2
Rp 1 2 6445.91
Cp 1 2 6.04p
Rs 1 N3 0.215
L1 N3 2 8.09u
.ends 4020_74437324100_10u 
*******
.subckt 4020_74437324150_15u  1 2
Rp 1 2 22764
Cp 1 2 5.34p
Rs 1 N3 0.325
L1 N3 2 13.18u
.ends 4020_74437324150_15u 
*******
.subckt 4020_74437324220_22u  1 2
Rp 1 2 11991.27
Cp 1 2 6.28p
Rs 1 N3 0.47
L1 N3 2 20.05u
.ends 4020_74437324220_22u 
*******
.subckt 4020_744373240010_0.1u  1 2
Rp 1 2 231.51
Cp 1 2 2.53p
Rs 1 N3 0.0032
L1 N3 2 0.092u
.ends 4020_744373240010_0.1u 
*******
.subckt 4020_744373240022_0.22u  1 2
Rp 1 2 339.47
Cp 1 2 3.64p
Rs 1 N3 0.0066
L1 N3 2 0.19u
.ends 4020_744373240022_0.22u 
*******
.subckt 4020_744373240033_0.33u  1 2
Rp 1 2 482.64
Cp 1 2 4.14p
Rs 1 N3 0.0078
L1 N3 2 0.3u
.ends 4020_744373240033_0.33u 
*******
.subckt 4020_744373240047_0.47u  1 2
Rp 1 2 614.49
Cp 1 2 4.59p
Rs 1 N3 0.0112
L1 N3 2 0.39u
.ends 4020_744373240047_0.47u 
*******
.subckt 4020_744373240056_0.56u  1 2
Rp 1 2 660.16
Cp 1 2 4.78p
Rs 1 N3 0.0135
L1 N3 2 0.51u
.ends 4020_744373240056_0.56u 
*******
.subckt 4020_744373240068_0.68u  1 2
Rp 1 2 1151.23
Cp 1 2 4.8226p
Rs 1 N3 0.016
L1 N3 2 0.63u
.ends 4020_744373240068_0.68u 
*******
.subckt 5020_74437334010_1u  1 2
Rp 1 2 2560.871340738
Cp 1 2 6.3479583446p
Rs 1 N3 0.0175
L1 N3 2 0.98u
.ends 5020_74437334010_1u 
*******
.subckt 5020_74437334012_1.2u  1 2
Rp 1 2 2938.105755004
Cp 1 2 5.8331555026p
Rs 1 N3 0.023
L1 N3 2 1.17u
.ends 5020_74437334012_1.2u 
*******
.subckt 5020_74437334015_1.5u  1 2
Rp 1 2 1600
Cp 1 2 13.5p
Rs 1 N3 0.0265
L1 N3 2 1.52u
.ends 5020_74437334015_1.5u 
*******
.subckt 5020_74437334022_2.2u  1 2
Rp 1 2 5165
Cp 1 2 5.925355369p
Rs 1 N3 0.042
L1 N3 2 2u
.ends 5020_74437334022_2.2u 
*******
.subckt 5020_74437334033_3.3u  1 2
Rp 1 2 7014.999879904
Cp 1 2 6.9257220898p
Rs 1 N3 0.066
L1 N3 2 3.04u
.ends 5020_74437334033_3.3u 
*******
.subckt 5020_74437334047_4.7u  1 2
Rp 1 2 9832.83582577
Cp 1 2 6.991567086p
Rs 1 N3 0.103
L1 N3 2 4.84u
.ends 5020_74437334047_4.7u 
*******
.subckt 5020_74437334056_5.6u  1 2
Rp 1 2 8004.185733344
Cp 1 2 9.3404220332p
Rs 1 N3 0.112
L1 N3 2 5.75u
.ends 5020_74437334056_5.6u 
*******
.subckt 5020_74437334068_6.8u  1 2
Rp 1 2 12363.72479874
Cp 1 2 9.0573395976p
Rs 1 N3 0.13
L1 N3 2 6.47u
.ends 5020_74437334068_6.8u 
*******
.subckt 5020_74437334082_8.2u  1 2
Rp 1 2 14406.34850544
Cp 1 2 6.8186289076p
Rs 1 N3 0.148
L1 N3 2 7.43u
.ends 5020_74437334082_8.2u 
*******
.subckt 5020_74437334100_10u  1 2
Rp 1 2 16863
Cp 1 2 8.51p
Rs 1 N3 0.18
L1 N3 2 10.32u
.ends 5020_74437334100_10u 
*******
.subckt 5020_744373340033_0.33u  1 2
Rp 1 2 9779.93165117333
Cp 1 2 6.94345698933333p
Rs 1 N3 0.0063
L1 N3 2 0.33u
.ends 5020_744373340033_0.33u 
*******
.subckt 5020_744373340047_0.47u  1 2
Rp 1 2 1116.67675146
Cp 1 2 6.6123463514p
Rs 1 N3 0.0073
L1 N3 2 0.44u
.ends 5020_744373340047_0.47u 
*******
.subckt 5020_744373340068_0.68u  1 2
Rp 1 2 1593.932714896
Cp 1 2 5.228244879p
Rs 1 N3 0.011
L1 N3 2 0.62u
.ends 5020_744373340068_0.68u 
*******
.subckt 5030_74437336010_1u  1 2
Rp 1 2 2437.684024608
Cp 1 2 7.0810090612p
Rs 1 N3 0.013
L1 N3 2 0.96u
.ends 5030_74437336010_1u 
*******
.subckt 5030_74437336012_1.2u  1 2
Rp 1 2 2220.61476690833
Cp 1 2 8.2230998956p
Rs 1 N3 0.014
L1 N3 2 1.26u
.ends 5030_74437336012_1.2u 
*******
.subckt 5030_74437336015_1.5u  1 2
Rp 1 2 3591.674613612
Cp 1 2 7.768760569p
Rs 1 N3 0.016
L1 N3 2 1.49u
.ends 5030_74437336015_1.5u 
*******
.subckt 5030_74437336022_2.2u  1 2
Rp 1 2 2670.312818732
Cp 1 2 7.4263445314p
Rs 1 N3 0.025
L1 N3 2 1.95u
.ends 5030_74437336022_2.2u 
*******
.subckt 5030_74437336033_3.3u  1 2
Rp 1 2 5773.34718188
Cp 1 2 9.579731907p
Rs 1 N3 0.032
L1 N3 2 3.29u
.ends 5030_74437336033_3.3u 
*******
.subckt 5030_74437336047_4.7u  1 2
Rp 1 2 6984.60185466
Cp 1 2 9.5379201058p
Rs 1 N3 0.05
L1 N3 2 4.35u
.ends 5030_74437336047_4.7u 
*******
.subckt 5030_74437336056_5.6u  1 2
Rp 1 2 8436.621935378
Cp 1 2 8.9830022734p
Rs 1 N3 0.055
L1 N3 2 5.7u
.ends 5030_74437336056_5.6u 
*******
.subckt 5030_74437336068_6.8u  1 2
Rp 1 2 3050
Cp 1 2 18.77p
Rs 1 N3 0.068
L1 N3 2 6.58u
.ends 5030_74437336068_6.8u 
*******
.subckt 5030_74437336100_10u  1 2
Rp 1 2 8904.428839494
Cp 1 2 9.050439242p
Rs 1 N3 0.11
L1 N3 2 10.44u
.ends 5030_74437336100_10u 
*******
.subckt 5030_744373360033_0.33u  1 2
Rp 1 2 484
Cp 1 2 11.45p
Rs 1 N3 0.0043
L1 N3 2 0.33u
.ends 5030_744373360033_0.33u 
*******
.subckt 5030_744373360047_0.47u  1 2
Rp 1 2 1270.694684518
Cp 1 2 5.7931935162p
Rs 1 N3 0.0064
L1 N3 2 0.46u
.ends 5030_744373360047_0.47u 
*******
.subckt 5030_744373360068_0.68u  1 2
Rp 1 2 1169.058072556
Cp 1 2 5.4791944186p
Rs 1 N3 0.01
L1 N3 2 0.59u
.ends 5030_744373360068_0.68u 
*******
.subckt 7030_74437346010_1u  1 2
Rp 1 2 1055.93
Cp 1 2 8.86p
Rs 1 N3 0.0083
L1 N3 2 1u
.ends 7030_74437346010_1u 
*******
.subckt 7030_74437346015_1.5u  1 2
Rp 1 2 1341.01
Cp 1 2 9.61p
Rs 1 N3 0.013
L1 N3 2 1.29u
.ends 7030_74437346015_1.5u 
*******
.subckt 7030_74437346018_1.8u  1 2
Rp 1 2 1489.8
Cp 1 2 11.46p
Rs 1 N3 0.014
L1 N3 2 1.69u
.ends 7030_74437346018_1.8u 
*******
.subckt 7030_74437346022_2.2u  1 2
Rp 1 2 1713.16
Cp 1 2 12.67p
Rs 1 N3 0.018
L1 N3 2 1.91u
.ends 7030_74437346022_2.2u 
*******
.subckt 7030_74437346025_2.5u  1 2
Rp 1 2 2127.67
Cp 1 2 12.13p
Rs 1 N3 0.02
L1 N3 2 2.4u
.ends 7030_74437346025_2.5u 
*******
.subckt 7030_74437346033_3.3u  1 2
Rp 1 2 3286.73
Cp 1 2 11.538p
Rs 1 N3 0.028
L1 N3 2 3.09u
.ends 7030_74437346033_3.3u 
*******
.subckt 7030_74437346047_4.7u  1 2
Rp 1 2 3661.93
Cp 1 2 12.75p
Rs 1 N3 0.037
L1 N3 2 4.22u
.ends 7030_74437346047_4.7u 
*******
.subckt 7030_74437346056_5.6u  1 2
Rp 1 2 3443.15
Cp 1 2 14.912p
Rs 1 N3 0.043
L1 N3 2 5.96u
.ends 7030_74437346056_5.6u 
*******
.subckt 7030_74437346068_6.8u  1 2
Rp 1 2 4377.18
Cp 1 2 12.16p
Rs 1 N3 0.054
L1 N3 2 6.19u
.ends 7030_74437346068_6.8u 
*******
.subckt 7030_74437346082_8.2u  1 2
Rp 1 2 3298.23
Cp 1 2 11.21p
Rs 1 N3 0.064
L1 N3 2 7.45u
.ends 7030_74437346082_8.2u 
*******
.subckt 7030_74437346100_10u  1 2
Rp 1 2 6696.59
Cp 1 2 13.59p
Rs 1 N3 0.075
L1 N3 2 8.42u
.ends 7030_74437346100_10u 
*******
.subckt 7030_74437346150_15u 1 2
Rp 1 2 10049
Cp 1 2 12.007p
Rs 1 N3 0.107
L1 N3 2 14.019u
.ends 7030_74437346150_15u
*******
.subckt 7030_74437346220_22u  1 2
Rp 1 2 9519.69
Cp 1 2 13.59p
Rs 1 N3 0.165
L1 N3 2 18.87u
.ends 7030_74437346220_22u 
*******
.subckt 7030_744373460022_0.22u  1 2
Rp 1 2 364.1
Cp 1 2 5.62p
Rs 1 N3 0.0021
L1 N3 2 0.2u
.ends 7030_744373460022_0.22u 
*******
.subckt 7030_744373460033_0.33u  1 2
Rp 1 2 478.45
Cp 1 2 5.67p
Rs 1 N3 0.0035
L1 N3 2 0.29u
.ends 7030_744373460033_0.33u 
*******
.subckt 7030_744373460047_0.47u  1 2
Rp 1 2 595.7
Cp 1 2 7.39p
Rs 1 N3 0.004
L1 N3 2 0.43u
.ends 7030_744373460047_0.47u 
*******
.subckt 7030_744373460068_0.68u  1 2
Rp 1 2 673.07
Cp 1 2 9.1p
Rs 1 N3 0.0048
L1 N3 2 0.54u
.ends 7030_744373460068_0.68u 
*******
.subckt 7030_744373460082_0.82u  1 2
Rp 1 2 875.76
Cp 1 2 9.4p
Rs 1 N3 0.0067
L1 N3 2 0.76u
.ends 7030_744373460082_0.82u 
*******
.subckt 7050_74437349010_1u  1 2
Rp 1 2 1144.82
Cp 1 2 9.89p
Rs 1 N3 0.0061
L1 N3 2 0.99u
.ends 7050_74437349010_1u 
*******
.subckt 7050_74437349012_1.2u  1 2
Rp 1 2 1314.53
Cp 1 2 10.42p
Rs 1 N3 0.0072
L1 N3 2 1.2u
.ends 7050_74437349012_1.2u 
*******
.subckt 7050_74437349015_1.5u  1 2
Rp 1 2 1285.43
Cp 1 2 14.07p
Rs 1 N3 0.0086
L1 N3 2 1.51u
.ends 7050_74437349015_1.5u 
*******
.subckt 7050_74437349022_2.2u  1 2
Rp 1 2 2074.35
Cp 1 2 12.82p
Rs 1 N3 0.0112
L1 N3 2 2.31u
.ends 7050_74437349022_2.2u 
*******
.subckt 7050_74437349033_3.3u  1 2
Rp 1 2 2798.93
Cp 1 2 12.21p
Rs 1 N3 0.019
L1 N3 2 3.11u
.ends 7050_74437349033_3.3u 
*******
.subckt 7050_74437349047_4.7u  1 2
Rp 1 2 3986.67
Cp 1 2 10.29p
Rs 1 N3 0.028
L1 N3 2 4.45u
.ends 7050_74437349047_4.7u 
*******
.subckt 7050_74437349056_5.6u  1 2
Rp 1 2 4945.14
Cp 1 2 13.22p
Rs 1 N3 0.044
L1 N3 2 6.31u
.ends 7050_74437349056_5.6u 
*******
.subckt 7050_74437349068_6.8u  1 2
Rp 1 2 5527.57
Cp 1 2 13.84p
Rs 1 N3 0.046
L1 N3 2 6.98u
.ends 7050_74437349068_6.8u 
*******
.subckt 7050_74437349082_8.2u  1 2
Rp 1 2 6412.43
Cp 1 2 14.82p
Rs 1 N3 0.056
L1 N3 2 7.88u
.ends 7050_74437349082_8.2u 
*******
.subckt 7050_74437349100_10u  1 2
Rp 1 2 8000
Cp 1 2 16p
Rs 1 N3 0.065
L1 N3 2 11.28u
.ends 7050_74437349100_10u 
*******
.subckt 7050_74437349150_15u  1 2
Rp 1 2 7092.51
Cp 1 2 15.05p
Rs 1 N3 0.081
L1 N3 2 14.76u
.ends 7050_74437349150_15u 
*******
.subckt 7050_74437349220_22u  1 2
Rp 1 2 11837.07
Cp 1 2 18.04p
Rs 1 N3 0.14
L1 N3 2 22.76u
.ends 7050_74437349220_22u 
*******
.subckt 7050_74437349330_33u  1 2
Rp 1 2 15573
Cp 1 2 13.208p
Rs 1 N3 0.173
L1 N3 2 35.22u
.ends 7050_74437349330_33u 
*******
.subckt 7050_74437349470_47u  1 2
Rp 1 2 32440
Cp 1 2 11.25p
Rs 1 N3 0.29
L1 N3 2 42.9u
.ends 7050_74437349470_47u 
*******
.subckt 7050_74437349560_56u  1 2
Rp 1 2 26898
Cp 1 2 12.58p
Rs 1 N3 0.342
L1 N3 2 59.42u
.ends 7050_74437349560_56u 
*******
.subckt 7050_74437349680_68u  1 2
Rp 1 2 18182
Cp 1 2 15.57p
Rs 1 N3 0.386
L1 N3 2 72.94u
.ends 7050_74437349680_68u 
*******
.subckt 7050_744373490047_0.47u  1 2
Rp 1 2 713.05
Cp 1 2 5.84p
Rs 1 N3 0.0035
L1 N3 2 0.45u
.ends 7050_744373490047_0.47u 
*******
.subckt 7050_744373490056_0.56u  1 2
Rp 1 2 681.13
Cp 1 2 7.03p
Rs 1 N3 0.0036
L1 N3 2 0.52u
.ends 7050_744373490056_0.56u 
*******
.subckt 7050_744373490068_0.68u  1 2
Rp 1 2 788.55
Cp 1 2 6.99p
Rs 1 N3 0.004
L1 N3 2 0.62u
.ends 7050_744373490068_0.68u 
*******
.subckt 7050_744373490082_0.82u  1 2
Rp 1 2 866.53
Cp 1 2 7.12p
Rs 1 N3 0.0046
L1 N3 2 0.72u
.ends 7050_744373490082_0.82u 
*******
.subckt 8030_74437356010_1u  1 2
Rp 1 2 1225.02497413
Cp 1 2 13.74399161p
Rs 1 N3 0.0051
L1 N3 2 0.92u
.ends 8030_74437356010_1u 
*******
.subckt 8030_74437356015_1.5u  1 2
Rp 1 2 1569.36944329
Cp 1 2 16.435199417p
Rs 1 N3 0.0083
L1 N3 2 1.6u
.ends 8030_74437356015_1.5u 
*******
.subckt 8030_74437356022_2.2u  1 2
Rp 1 2 1989.16375073
Cp 1 2 18.489074561p
Rs 1 N3 0.0136
L1 N3 2 2.5u
.ends 8030_74437356022_2.2u 
*******
.subckt 8030_74437356033_3.3u  1 2
Rp 1 2 2469.55214706667
Cp 1 2 19.7843439316667p
Rs 1 N3 0.0188
L1 N3 2 3.56u
.ends 8030_74437356033_3.3u 
*******
.subckt 8030_74437356047_4.7u  1 2
Rp 1 2 1532.12191441
Cp 1 2 21.911597874p
Rs 1 N3 0.0266
L1 N3 2 4.2u
.ends 8030_74437356047_4.7u 
*******
.subckt 8030_74437356068_6.8u  1 2
Rp 1 2 2112.78616687
Cp 1 2 20.477571059p
Rs 1 N3 0.0355
L1 N3 2 6.1u
.ends 8030_74437356068_6.8u 
*******
.subckt 8030_74437356082_8.2u  1 2
Rp 1 2 2401.7535144
Cp 1 2 22.791773101p
Rs 1 N3 0.0564
L1 N3 2 8.98u
.ends 8030_74437356082_8.2u 
*******
.subckt 8030_74437356100_10u  1 2
Rp 1 2 2434.5525673
Cp 1 2 25.978385807p
Rs 1 N3 0.061
L1 N3 2 10.59u
.ends 8030_74437356100_10u 
*******
.subckt 8030_744373560022_0.22u  1 2
Rp 1 2 335.009326058
Cp 1 2 9.525394418p
Rs 1 N3 0.00147
L1 N3 2 0.2u
.ends 8030_744373560022_0.22u 
*******
.subckt 8030_744373560033_0.33u  1 2
Rp 1 2 620.655456145
Cp 1 2 9.576544239p
Rs 1 N3 0.00206
L1 N3 2 0.33u
.ends 8030_744373560033_0.33u 
*******
.subckt 8030_744373560047_0.47u  1 2
Rp 1 2 628.753910793
Cp 1 2 11.257388855p
Rs 1 N3 0.00235
L1 N3 2 0.42u
.ends 8030_744373560047_0.47u 
*******
.subckt 8030_744373560068_0.68u  1 2
Rp 1 2 882.559693359
Cp 1 2 12.77945307p
Rs 1 N3 0.00365
L1 N3 2 0.69u
.ends 8030_744373560068_0.68u 
*******
.subckt 8030_744373560082_0.82u  1 2
Rp 1 2 1004.98958848
Cp 1 2 12.256703154p
Rs 1 N3 0.0042
L1 N3 2 0.75u
.ends 8030_744373560082_0.82u 
*******
.subckt 8040_74437358010_1u  1 2
Rp 1 2 1309.95123894
Cp 1 2 14.8796442454p
Rs 1 N3 0.00365
L1 N3 2 0.97u
.ends 8040_74437358010_1u 
*******
.subckt 8040_74437358022_2.2u  1 2
Rp 1 2 1655.969312838
Cp 1 2 15.2109156398p
Rs 1 N3 0.0087
L1 N3 2 2.07u
.ends 8040_74437358022_2.2u 
*******
.subckt 8040_74437358033_3.3u  1 2
Rp 1 2 1504.6
Cp 1 2 19.8812p
Rs 1 N3 0.01235
L1 N3 2 3.85u
.ends 8040_74437358033_3.3u 
*******
.subckt 8040_74437358047_4.7u  1 2
Rp 1 2 4606.353956504
Cp 1 2 17.1496262976p
Rs 1 N3 0.0197
L1 N3 2 5.4u
.ends 8040_74437358047_4.7u 
*******
.subckt 8040_74437358068_6.8u  1 2
Rp 1 2 2785.289422032
Cp 1 2 25.3812020296p
Rs 1 N3 0.0292
L1 N3 2 6.64u
.ends 8040_74437358068_6.8u 
*******
.subckt 8040_74437358082_8.2u  1 2
Rp 1 2 9109.407410496
Cp 1 2 24.7673114866p
Rs 1 N3 0.0411
L1 N3 2 9.49u
.ends 8040_74437358082_8.2u 
*******
.subckt 8040_74437358100_10u  1 2
Rp 1 2 2613.576862176
Cp 1 2 29.3485071434p
Rs 1 N3 0.0481
L1 N3 2 10.7u
.ends 8040_74437358100_10u 
*******
.subckt 8040_744373580022_0.22u  1 2
Rp 1 2 501.3260830762
Cp 1 2 7.049576596p
Rs 1 N3 0.00087
L1 N3 2 0.19u
.ends 8040_744373580022_0.22u 
*******
.subckt 8040_744373580033_0.33u  1 2
Rp 1 2 718.767385631
Cp 1 2 8.4782375374p
Rs 1 N3 0.00145
L1 N3 2 0.34u
.ends 8040_744373580033_0.33u 
*******
.subckt 8040_744373580047_0.47u  1 2
Rp 1 2 783.9580966398
Cp 1 2 9.6095127766p
Rs 1 N3 0.00168
L1 N3 2 0.45u
.ends 8040_744373580047_0.47u 
*******
.subckt 8040_744373580068_0.68u  1 2
Rp 1 2 795.4562492636
Cp 1 2 16.5237360048p
Rs 1 N3 0.00275
L1 N3 2 0.73u
.ends 8040_744373580068_0.68u 
*******
.subckt 8040_744373580082_0.82u  1 2
Rp 1 2 902.7579230984
Cp 1 2 13.4922532316p
Rs 1 N3 0.00295
L1 N3 2 0.72u
.ends 8040_744373580082_0.82u 
*******
