**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Auxiliary Gate Drive Transformer
* Matchcode:              WE-AGDT
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Toby      
* Date and Time:          2022-06-29
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************		
.subckt	750317893		1  3  2  4  8  5		
.param RxLkg=875.14ohm					
.param Leakage=0.328uh					
Rlkg	1	1a	{RxLkg*2}		
L_Lkg	1	1a	{Leakage*2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg*2}		
L_Lkg2	2	2a	{Leakage*2}	Rser=0.01mohm	
Lpri1	1a	3	17.672uH	Rser=166mohm	
Lpri2	2a	4	17.672uH	Rser=166mohm	
Lsec1	8	5	72uH	Rser=395mohm	
K Lpri1 Lpri2   Lsec1        1					
.param Cprm1=9.755pf					
.param Cprm2=9.755pf					
.param Rdmp1=48026.1ohm					
.param Rdmp2=48026.1ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Cpri2	2	4	{Cprm2}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rdmp2	2	4	{Rdmp2}		
Rg3	1	0	20meg		
Rg4	2	0	20meg		
Rg7	3	0	20meg		
Rg8	4	0	20meg		
Rg11	8	0	20meg		
Rg19	5	0	20meg		
.ends		


.subckt	750317894		1  4  8  5  7  6		
.param RxLkg=1097.35ohm					
.param Leakage=0.255uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	4	17.745uH	Rser=85mohm	
Lsec1	8	5	43.556uH	Rser=260mohm	
Lsec2	7	6	3.556uH	Rser=85mohm	
K Lpri1    Lsec1 Lsec2       1					
.param Cprm1=7.5pf					
.param Rdmp1=77459.69ohm					
Cpri1	1	4	{Cprm1}	Rser=10mohm	
Rdmp1	1	4	{Rdmp1}		
Rg3	1	0	20meg		
Rg7	4	0	20meg		
Rg11	8	0	20meg		
Rg12	7	0	20meg		
Rg19	5	0	20meg		
Rg20	6	0	20meg		
.ends	


.subckt	750318114		1  3  2  4  8  6		
.param RxLkg=1249.42ohm					
.param Leakage=0.285uh					
Rlkg	1	1a	{RxLkg*2}		
L_Lkg	1	1a	{Leakage*2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg*2}		
L_Lkg2	2	2a	{Leakage*2}	Rser=0.01mohm	
Lpri1	1a	3	5.715uH	Rser=120mohm	
Lpri2	2a	4	5.715uH	Rser=120mohm	
Lsec1	8	6	24uH	Rser=285mohm	
K Lpri1 Lpri2   Lsec1        1					
.param Cprm1=10.84pf					
.param Cprm2=10.84pf					
.param Rdmp1=26303.65ohm					
.param Rdmp2=26303.65ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Cpri2	2	4	{Cprm2}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rdmp2	2	4	{Rdmp2}		
Rg3	1	0	20meg		
Rg4	2	0	20meg		
Rg7	3	0	20meg		
Rg8	4	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends	

		
.subckt	750318131		1  3  2  4  8  6  7  5		
.param RxLkg=1517.91ohm					
.param Leakage=0.27uh					
Rlkg	1	1a	{RxLkg*2}		
L_Lkg	1	1a	{Leakage*2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg*2}		
L_Lkg2	2	2a	{Leakage*2}	Rser=0.01mohm	
Lpri1	1a	3	6.73uH	Rser=94mohm	
Lpri2	2a	4	6.73uH	Rser=94mohm	
Lsec1	8	6	16.938uH	Rser=205mohm	
Lsec2	7	5	1.383uH	Rser=71mohm	
K Lpri1 Lpri2   Lsec1 Lsec2       1					
.param Cprm1=5.65pf					
.param Cprm2=5.65pf					
.param Rdmp1=39353.16ohm					
.param Rdmp2=39353.16ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Cpri2	2	4	{Cprm2}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rdmp2	2	4	{Rdmp2}		
Rg3	1	0	20meg		
Rg4	2	0	20meg		
Rg7	3	0	20meg		
Rg8	4	0	20meg		
Rg11	8	0	20meg		
Rg12	7	0	20meg		
Rg19	6	0	20meg		
Rg20	5	0	20meg		
.ends	
		

.subckt	750318207		1  4  8  5		
.param RxLkg=1822.36ohm					
.param Leakage=0.539uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	4	26.461uH	Rser=240mohm	
Lsec1	8	5	38.88uH	Rser=353mohm	
K Lpri1    Lsec1        1					
.param Cprm1=8.1pf					
.param Rdmp1=91287.02ohm					
Cpri1	1	4	{Cprm1}	Rser=10mohm	
Rdmp1	1	4	{Rdmp1}		
Rg3	1	0	20meg		
Rg7	4	0	20meg		
Rg11	8	0	20meg		
Rg19	5	0	20meg		
.ends					
		
	
.subckt	750318208		1  4  8  5  7  6		
.param RxLkg=1748.22ohm					
.param Leakage=0.325uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	4	26.675uH	Rser=155mohm	
Lsec1	8	5	27uH	Rser=250mohm	
Lsec2	7	6	2.204uH	Rser=85mohm	
K Lpri1    Lsec1 Lsec2       1					
.param Cprm1=3.2pf					
.param Rdmp1=145236.83ohm					
Cpri1	1	4	{Cprm1}	Rser=10mohm	
Rdmp1	1	4	{Rdmp1}		
Rg3	1	0	20meg		
Rg7	4	0	20meg		
Rg11	8	0	20meg		
Rg12	7	0	20meg		
Rg19	5	0	20meg		
Rg20	6	0	20meg		
.ends		


.subckt	750318616		1  3  2  4  8  5		
.param RxLkg=585.54ohm					
.param Leakage=0.12uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	9.88uH	Rser=50mohm	
Laux1	2	4	6.944uH	Rser=104mohm	
Lsec1	8	5	27.778uH	Rser=260mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=10.5pf					
.param Rdmp1=48795.03ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	2	0	20meg		
Rg7	3	0	20meg		
Rg9	4	0	20meg		
Rg11	8	0	20meg		
Rg19	5	0	20meg		
.ends	



.subckt	750319077		2  1  4  3  5  6  7  8		
.param RxLkg=568.63ohm					
.param Leakage=0.39uh					
Rlkg	2	2a	{RxLkg}		
L_Lkg	2	2a	{Leakage}	Rser=0.01mohm	
Lpri1	2a	1	41.61uH	Rser=195mohm	
Laux1	4	3	10.5uH	Rser=132mohm	
Lsec1	5	6	85.714uH	Rser=1300mohm	
Lsec2	7	6	21.429uH	Rser=700mohm	
Lsec3	6	8	21.429uH	Rser=700mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=28pf					
.param Rdmp1=61237.34ohm					
Cpri1	2	1	{Cprm1}	Rser=10mohm	
Rdmp1	2	1	{Rdmp1}		
Rg3	2	0	20meg		
Rg5	4	0	20meg		
Rg7	1	0	20meg		
Rg9	3	0	20meg		
Rg11	5	0	20meg		
Rg12	7	0	20meg		
Rg19	6	0	20meg			
Rg21	8	0	20meg		
.ends					
			

.subckt	750319177		1  3  8  6		
.param RxLkg=1513.83ohm					
.param Leakage=0.55uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	29.45uH	Rser=45mohm	
Lsec1	8	6	83.333uH	Rser=115mohm	
K Lpri1    Lsec1        1					
.param Cprm1=11pf					
.param Rdmp1=82572.36ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg7	3	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends					
							

.subckt	750319282		2  1  4  3  5  6  7  8		
.param RxLkg=586.95ohm					
.param Leakage=0.65uh					
Rlkg	2	2a	{RxLkg}		
L_Lkg	2	2a	{Leakage}	Rser=0.01mohm	
Lpri1	2a	1	41.35uH	Rser=215mohm	
Laux1	4	3	17.357uH	Rser=196mohm	
Lsec1	5	6	262.5uH	Rser=2400mohm	
Lsec2	6	8	17.357uH	Rser=660mohm	
Lsec3	7	6	17.357uH	Rser=660mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=73pf					
.param Rdmp1=37925.76ohm					
Cpri1	2	1	{Cprm1}	Rser=10mohm	
Rdmp1	2	1	{Rdmp1}		
Rg3	2	0	20meg		
Rg5	4	0	20meg		
Rg7	1	0	20meg		
Rg9	3	0	20meg		
Rg11	5	0	20meg		
Rg13	7	0	20meg		
Rg19	6	0	20meg		
Rg20	8	0	20meg			
.ends					
		

.subckt	750319331		1  3  8  6		
.param RxLkg=2970.44ohm					
.param Leakage=1.5uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	73.5uH	Rser=85mohm	
Lsec1	8	6	75uH	Rser=85mohm	
K Lpri1    Lsec1        1					
.param Cprm1=8.5pf					
.param Rdmp1=148522.25ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg7	3	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends								
	

.subckt	750319496		1  3  8  6  7  5		
.param RxLkg=1192.28ohm					
.param Leakage=0.275uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	6.725uH	Rser=42mohm	
Lsec1	8	6	28uH	Rser=370mohm	
Lsec2	7	5	2.16uH	Rser=115mohm	
K Lpri1    Lsec1 Lsec2       1					
.param Cprm1=19pf					
.param Rdmp1=30348.84ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg7	3	0	20meg		
Rg11	8	0	20meg		
Rg12	7	0	20meg		
Rg19	6	0	20meg		
Rg20	5	0	20meg		
.ends					


.subckt	750319497		1  3  8  6  7  5		
.param RxLkg=1122.95ohm					
.param Leakage=0.245uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	6.755uH	Rser=42mohm	
Lsec1	8	6	24.975uH	Rser=350mohm	
Lsec2	7	5	1.383uH	Rser=95mohm	
K Lpri1    Lsec1 Lsec2       1					
.param Cprm1=17pf					
.param Rdmp1=32084.43ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg7	3	0	20meg		
Rg11	8	0	20meg		
Rg12	7	0	20meg		
Rg19	6	0	20meg		
Rg20	5	0	20meg		
.ends					
		

.subckt	750319565		1  3  8  6		
.param RxLkg=1562.5ohm					
.param Leakage=2.5uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	253.5uH	Rser=275mohm	
Lsec1	8	6	1024uH	Rser=345mohm	
K Lpri1    Lsec1        1					
.param Cprm1=25pf					
.param Rdmp1=160000.26ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg7	3	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends