**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  Aluminum Electrolytic Capacitors
* Matchcode:              WCAP-AIG8
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/21/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 861010784009_3.3mF 1 2
Rser 1 3 0.04072
Lser 2 4 2.1779506405E-08
C1 3 4 0.0033
Rpar 3 4 15151.5151515152
.ends 861010784009_3.3mF
*******
.subckt 861010786015_4.7mF 1 2
Rser 1 3 0.037283
Lser 2 4 1.9842938336E-08
C1 3 4 0.0047
Rpar 3 4 10638.2978723404
.ends 861010786015_4.7mF
*******
.subckt 861010786021_6.8mF 1 2
Rser 1 3 0.037173
Lser 2 4 1.9088268647E-08
C1 3 4 0.0068
Rpar 3 4 7352.94117647059
.ends 861010786021_6.8mF
*******
.subckt 861011084009_470uF 1 2
Rser 1 3 0.1485
Lser 2 4 1.6657293561E-08
C1 3 4 0.00047
Rpar 3 4 106382.978723404
.ends 861011084009_470uF
*******
.subckt 861011084015_680uF 1 2
Rser 1 3 0.12221
Lser 2 4 1.6423797781E-08
C1 3 4 0.00068
Rpar 3 4 73529.4117647059
.ends 861011084015_680uF
*******
.subckt 861011086027_1.5mF 1 2
Rser 1 3 0.060055
Lser 2 4 1.7054937341E-08
C1 3 4 0.0015
Rpar 3 4 33333.3333333333
.ends 861011086027_1.5mF
*******
.subckt 861011384014_220uF 1 2
Rser 1 3 0.31844
Lser 2 4 1.4863233484E-08
C1 3 4 0.00022
Rpar 3 4 227272.727272727
.ends 861011384014_220uF
*******
.subckt 861011385023_330uF 1 2
Rser 1 3 0.22242
Lser 2 4 1.2037845668E-08
C1 3 4 0.00033
Rpar 3 4 151515.151515152
.ends 861011385023_330uF
*******
.subckt 861011386030_470uF 1 2
Rser 1 3 0.17265
Lser 2 4 1.3520559628E-08
C1 3 4 0.00047
Rpar 3 4 106382.978723404
.ends 861011386030_470uF
*******
.subckt 861011483001_47uF 1 2
Rser 1 3 0.592
Lser 2 4 1.3511713379E-08
C1 3 4 0.000047
Rpar 3 4 1063829.78723404
.ends 861011483001_47uF
*******
.subckt 861011483002_68uF 1 2
Rser 1 3 0.592
Lser 2 4 1.3027728829E-08
C1 3 4 0.000068
Rpar 3 4 735294.117647059
.ends 861011483002_68uF
*******
.subckt 861011483003_82uF 1 2
Rser 1 3 0.298
Lser 2 4 1.3853014923E-08
C1 3 4 0.000082
Rpar 3 4 609756.097560976
.ends 861011483003_82uF
*******
.subckt 861011483004_100uF 1 2
Rser 1 3 0.26
Lser 2 4 1.2322764467E-08
C1 3 4 0.0001
Rpar 3 4 500000
.ends 861011483004_100uF
*******
.subckt 861011483005_120uF 1 2
Rser 1 3 0.213
Lser 2 4 1.3381590937E-08
C1 3 4 0.00012
Rpar 3 4 416666.666666667
.ends 861011483005_120uF
*******
.subckt 861011483006_150uF 1 2
Rser 1 3 0.188
Lser 2 4 1.3236124722E-08
C1 3 4 0.00015
Rpar 3 4 333333.333333333
.ends 861011483006_150uF
*******
.subckt 861011483007_180uF 1 2
Rser 1 3 0.163
Lser 2 4 1.2671116928E-08
C1 3 4 0.00018
Rpar 3 4 277777.777777778
.ends 861011483007_180uF
*******
.subckt 861011484008_82uF 1 2
Rser 1 3 0.346
Lser 2 4 1.5008879464E-08
C1 3 4 0.000082
Rpar 3 4 609756.097560976
.ends 861011484008_82uF
*******
.subckt 861011484009_100uF 1 2
Rser 1 3 0.262
Lser 2 4 1.90248154153584E-08
C1 3 4 0.0001
Rpar 3 4 500000
.ends 861011484009_100uF
*******
.subckt 861011484010_120uF 1 2
Rser 1 3 0.246
Lser 2 4 1.85213187898072E-08
C1 3 4 0.00012
Rpar 3 4 416666.666666667
.ends 861011484010_120uF
*******
.subckt 861011484011_150uF 1 2
Rser 1 3 0.183
Lser 2 4 1.3944336044E-08
C1 3 4 0.00015
Rpar 3 4 333333.333333333
.ends 861011484011_150uF
*******
.subckt 861011484012_180uF 1 2
Rser 1 3 0.152
Lser 2 4 1.3599919566E-08
C1 3 4 0.00018
Rpar 3 4 277777.777777778
.ends 861011484012_180uF
*******
.subckt 861011484013_220uF 1 2
Rser 1 3 0.127
Lser 2 4 1.35170052E-08
C1 3 4 0.00022
Rpar 3 4 227272.727272727
.ends 861011484013_220uF
*******
.subckt S861011784003_1.1mF 1 2
Rser 1 3 0.067
Lser 2 4 0.000000008
C1 3 4 0.0011
Rpar 3 4 89887.6404494382
.ends S861011784003_1.1mF
*******
.subckt 861011485014_150uF 1 2
Rser 1 3 0.205
Lser 2 4 2.45036491425324E-08
C1 3 4 0.00015
Rpar 3 4 333333.333333333
.ends 861011485014_150uF
*******
.subckt 861011485015_180uF 1 2
Rser 1 3 0.169
Lser 2 4 1.457289665E-08
C1 3 4 0.00018
Rpar 3 4 277777.777777778
.ends 861011485015_180uF
*******
.subckt 861011485016_220uF 1 2
Rser 1 3 0.148
Lser 2 4 2.47351457940872E-08
C1 3 4 0.00022
Rpar 3 4 227272.727272727
.ends 861011485016_220uF
*******
.subckt 861011485017_270uF 1 2
Rser 1 3 0.136
Lser 2 4 2.51911472421803E-08
C1 3 4 0.00027
Rpar 3 4 185185.185185185
.ends 861011485017_270uF
*******
.subckt 861011485018_330uF 1 2
Rser 1 3 0.121
Lser 2 4 2.61270674037942E-08
C1 3 4 0.00033
Rpar 3 4 151515.151515152
.ends 861011485018_330uF
*******
.subckt 861011485019_390uF 1 2
Rser 1 3 0.121
Lser 2 4 2.60587299530843E-08
C1 3 4 0.00039
Rpar 3 4 128205.128205128
.ends 861011485019_390uF
*******
.subckt 861011486020_220uF 1 2
Rser 1 3 0.31445
Lser 2 4 1.5829460581E-08
C1 3 4 0.00022
Rpar 3 4 227272.727272727
.ends 861011486020_220uF
*******
.subckt 861011486021_270uF 1 2
Rser 1 3 0.151
Lser 2 4 2.71212258520702E-08
C1 3 4 0.00027
Rpar 3 4 185185.185185185
.ends 861011486021_270uF
*******
.subckt 861011486022_330uF 1 2
Rser 1 3 0.104
Lser 2 4 9.09014270834679E-09
C1 3 4 0.00033
Rpar 3 4 151515.151515152
.ends 861011486022_330uF
*******
.subckt 861011486023_390uF 1 2
Rser 1 3 0.101
Lser 2 4 2.31407416896361E-08
C1 3 4 0.00039
Rpar 3 4 128205.128205128
.ends 861011486023_390uF
*******
.subckt 861011486024_470uF 1 2
Rser 1 3 0.076
Lser 2 4 9.10992922174604E-09
C1 3 4 0.00047
Rpar 3 4 106382.978723404
.ends 861011486024_470uF
*******
.subckt 861011487025_390uF 1 2
Rser 1 3 0.084
Lser 2 4 1.02705515973701E-08
C1 3 4 0.00039
Rpar 3 4 128205.128205128
.ends 861011487025_390uF
*******
.subckt 861011487026_470uF 1 2
Rser 1 3 0.082
Lser 2 4 1.0143049562128E-08
C1 3 4 0.00047
Rpar 3 4 106382.978723404
.ends 861011487026_470uF
*******
.subckt 861011487027_560uF 1 2
Rser 1 3 0.063
Lser 2 4 9.81318509955244E-09
C1 3 4 0.00056
Rpar 3 4 89285.7142857143
.ends 861011487027_560uF
*******
