**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Power Molded Chip Inductor
* Matchcode:              WE-PMCI 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0603_74479262147_0.47u 1 2
Rp 1 2 1100
Cp 1 2 1.7p
Rs 1 N3 0.087
L1 N3 2 0.47u
.ends 0603_74479262147_0.47u
*******
.subckt 0603_74479262210_1u 1 2
Rp 1 2 1900
Cp 1 2 2.8p
Rs 1 N3 0.17
L1 N3 2 1u
.ends 0603_74479262210_1u
*******
.subckt 0805_74479275147_0.47u 1 2
Rp 1 2 920
Cp 1 2 2.45p
Rs 1 N3 0.038
L1 N3 2 0.47u
.ends 0805_74479275147_0.47u
*******
.subckt 0805_74479275210_1u 1 2
Rp 1 2 1700
Cp 1 2 3.5p
Rs 1 N3 0.069
L1 N3 2 1u
.ends 0805_74479275210_1u
*******
.subckt 0805_74479275222_2.2u 1 2
Rp 1 2 2000
Cp 1 2 3.9p
Rs 1 N3 0.166
L1 N3 2 2.2u
.ends 0805_74479275222_2.2u
*******
.subckt 0806_74479276124_0.24u 1 2
Rp 1 2 600
Cp 1 2 2.4p
Rs 1 N3 0.019
L1 N3 2 0.24u
.ends 0806_74479276124_0.24u
*******
.subckt 0806_74479276147_0.47u 1 2
Rp 1 2 850
Cp 1 2 3p
Rs 1 N3 0.034
L1 N3 2 0.47u
.ends 0806_74479276147_0.47u
*******
.subckt 0806_74479276147C_0.47u 1 2
Rp 1 2 1000
Cp 1 2 3.3p
Rs 1 N3 0.033
L1 N3 2 0.47u
.ends 0806_74479276147C_0.47u
*******
.subckt 0806_74479276168_0.68u 1 2
Rp 1 2 1400
Cp 1 2 3p
Rs 1 N3 0.045
L1 N3 2 0.68u
.ends 0806_74479276168_0.68u
*******
.subckt 0806_74479276210_1u 1 2
Rp 1 2 1800
Cp 1 2 5p
Rs 1 N3 0.065
L1 N3 2 1u
.ends 0806_74479276210_1u
*******
.subckt 0806_74479276210C_1u 1 2
Rp 1 2 1500
Cp 1 2 4p
Rs 1 N3 0.053
L1 N3 2 1u
.ends 0806_74479276210C_1u
*******
.subckt 0806_74479276222_2.2u 1 2
Rp 1 2 3700
Cp 1 2 6p
Rs 1 N3 0.135
L1 N3 2 2.2u
.ends 0806_74479276222_2.2u
*******
.subckt 0806_74479276222C_2.2u 1 2
Rp 1 2 2500
Cp 1 2 4.5p
Rs 1 N3 0.112
L1 N3 2 2.2u
.ends 0806_74479276222C_2.2u
*******
.subckt 1008_74479287147_0.47u 1 2
Rp 1 2 1000
Cp 1 2 4p
Rs 1 N3 0.025
L1 N3 2 0.47u
.ends 1008_74479287147_0.47u
*******
.subckt 1008_74479287210_1u 1 2
Rp 1 2 1800
Cp 1 2 5p
Rs 1 N3 0.055
L1 N3 2 1u
.ends 1008_74479287210_1u
*******
.subckt 1008_74479287222_2.2u 1 2
Rp 1 2 3700
Cp 1 2 6p
Rs 1 N3 0.132
L1 N3 2 2.2u
.ends 1008_74479287222_2.2u
*******
.subckt 1008_74479288147_0.47u 1 2
Rp 1 2 1200
Cp 1 2 2p
Rs 1 N3 0.028
L1 N3 2 0.47u
.ends 1008_74479288147_0.47u
*******
.subckt 1008_74479288210_1u 1 2
Rp 1 2 1900
Cp 1 2 5.7p
Rs 1 N3 0.04
L1 N3 2 1u
.ends 1008_74479288210_1u
*******
.subckt 1008_74479288222_2.2u 1 2
Rp 1 2 3400
Cp 1 2 6.8p
Rs 1 N3 0.09
L1 N3 2 2.2u
.ends 1008_74479288222_2.2u
*******
.subckt 1008HS_74479288215_1.5u 1 2
Rp 1 2 2282
Cp 1 2 6.299p
Rs 1 N3 0.056
L1 N3 2 1.436u
.ends 1008HS_74479288215_1.5u
*******
.subckt 1210_74479298147_0.47u 1 2
Rp 1 2 920
Cp 1 2 5.1p
Rs 1 N3 0.028
L1 N3 2 0.47u
.ends 1210_74479298147_0.47u
*******
.subckt 1210_74479298210_1u 1 2
Rp 1 2 2200
Cp 1 2 5.3p
Rs 1 N3 0.045
L1 N3 2 1u
.ends 1210_74479298210_1u
*******
.subckt 1210_74479298222_2.2u 1 2
Rp 1 2 3600
Cp 1 2 7p
Rs 1 N3 0.096
L1 N3 2 2.2u
.ends 1210_74479298222_2.2u
*******
.subckt 1210_74479299147_0.47u 1 2
Rp 1 2 1000
Cp 1 2 4.8p
Rs 1 N3 0.025
L1 N3 2 0.47u
.ends 1210_74479299147_0.47u
*******
.subckt 1210_74479299210_1u 1 2
Rp 1 2 1700
Cp 1 2 6p
Rs 1 N3 0.038
L1 N3 2 1u
.ends 1210_74479299210_1u
*******
.subckt 1210_74479299222_2.2u 1 2
Rp 1 2 4000
Cp 1 2 7p
Rs 1 N3 0.085
L1 N3 2 2.2u
.ends 1210_74479299222_2.2u
*******
.subckt 1210HS_74479290125_0.25u 1 2
Rp 1 2 627.28
Cp 1 2 3.06p
Rs 1 N3 0.01
L1 N3 2 0.238u
.ends 1210HS_74479290125_0.25u
*******
