**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  Power over Ethernet Transformer
* Matchcode:              WE-PoE
* Library Type:           LTspice
* Version:                rev23b
* Created/modified by:    Roberta      
* Date and Time:          2023-03-07
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************	
* Copyright(C) 2023 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************
************ WE-PoE **************
.subckt	750315422		2  3  1  4  5  6  11  7		
.param RxLkg=154.84ohm					
.param Leakage=0.16uh					
Rlkg	2	2a	{RxLkg*2}		
L_Lkg	2	2a	{Leakage*2}	Rser=0.01mohm	
Rlkg2	1	1a	{RxLkg*2}		
L_Lkg2	1	1a	{Leakage*2}	Rser=0.01mohm	
Lpri1	2a	3	8.84uH	Rser=23mohm	
Lpri2	1a	4	8.84uH	Rser=27mohm	
Laux1	5	6	9uH	Rser=385mohm	
Lsec1	11	7	11.391uH	Rser=14mohm	
K Lpri1 Lpri2 Laux1  Lsec1        1					
.param Cprm1=148.3pf					
.param Cprm2=148.3pf					
.param Rdmp1=8709.74ohm					
.param Rdmp2=8709.74ohm					
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Cpri2	1	4	{Cprm2}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}		
Rdmp2	1	4	{Rdmp2}		
Rg3	2	0	20meg		
Rg4	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg8	4	0	20meg		
Rg9	6	0	20meg		
Rg11	11	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750313109		4  3  2  1  5  7  6  8		
.param RxLkg=3015.11ohm					
.param Leakage=0.8uh					
Rlkg	4	4a	{RxLkg}		
L_Lkg	4	4a	{Leakage}	Rser=0.01mohm	
Lpri1	4a	3	43.2uH	Rser=305mohm	
Laux1	2	1	17.188uH	Rser=438mohm	
Lsec1	5	7	2.75uH	Rser=40mohm	
Lsec2	6	8	2.75uH	Rser=40mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=4pf					
.param Rdmp1=165831.31ohm					
Cpri1	4	3	{Cprm1}	Rser=10mohm	
Rdmp1	4	3	{Rdmp1}		
Rg3	4	0	20meg		
Rg5	2	0	20meg		
Rg7	3	0	20meg		
Rg9	1	0	20meg		
Rg11	5	0	20meg		
Rg12	6	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
.ends					

.subckt	750344488		3  1  5  4  9  6		
.param RxLkg=255.83ohm					
.param Leakage=0.158uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	13.842uH	Rser=18mohm	
Laux1	5	4	7.875uH	Rser=126mohm	
Lsec1	9	6	7.875uH	Rser=13mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=68.11pf					
.param Rdmp1=22668.83ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	5	0	20meg		
Rg7	1	0	20meg		
Rg9	4	0	20meg		
Rg11	9	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt	750317123		2  1  3  4  6  7		
.param RxLkg=417.39ohm					
.param Leakage=0.6uh					
Rlkg	2	2a	{RxLkg}		
L_Lkg	2	2a	{Leakage}	Rser=0.01mohm	
Lpri1	2a	1	81.4uH	Rser=88mohm	
Laux1	3	4	7.38uH	Rser=56mohm	
Lsec1	6	7	13.12uH	Rser=16mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=63pf					
.param Rdmp1=57043.75ohm					
Cpri1	2	1	{Cprm1}	Rser=10mohm	
Rdmp1	2	1	{Rdmp1}		
Rg3	2	0	20meg		
Rg5	3	0	20meg		
Rg7	1	0	20meg		
Rg9	4	0	20meg		
Rg11	6	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310019		3  4  2  1  6  8  5  7		
.param RxLkg=4526.61ohm					
.param Leakage=4.5uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	305.5uH	Rser=1600mohm	
Laux1	2	1	576.446uH	Rser=2600mohm	
Lsec1	6	8	40.992uH	Rser=77.8mohm	
Lsec2	5	7	40.992uH	Rser=78.6mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=7.97pf					
.param Rdmp1=311832.98ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	6	0	20meg		
Rg12	5	0	20meg		
Rg19	8	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	750310018		3  4  2  1  5  7		
.param RxLkg=4601.31ohm					
.param Leakage=6.75uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	493.25uH	Rser=1570mohm	
Laux1	2	1	21.701uH	Rser=190mohm	
Lsec1	5	7	3.472uH	Rser=10mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=10.76pf					
.param Rdmp1=340837.67ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	5	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310022		3  4  2  1  5  7		
.param RxLkg=3999.97ohm					
.param Leakage=7.5uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	513.5uH	Rser=1600mohm	
Laux1	2	1	21.699uH	Rser=200mohm	
Lsec1	5	7	42.531uH	Rser=90mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=16.87pf					
.param Rdmp1=277864.58ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	5	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310020		3  4  2  1  5  7		
.param RxLkg=2940.26ohm					
.param Leakage=5.42uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	494.58uH	Rser=1620mohm	
Laux1	2	1	21.701uH	Rser=180mohm	
Lsec1	5	7	7.813uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=16.99pf					
.param Rdmp1=271241.97ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	5	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750314782		5  4  3  2  1  6  10  7  9		
.param RxLkg=470.46ohm					
.param Leakage=0.3uh					
Rlkg	5	5a	{RxLkg/2}		
L_Lkg	5	5a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	4	4a	{RxLkg/2}		
L_Lkg2	4	4a	{Leakage/2}	Rser=0.01mohm	
Lpri1	5a	4	9.1uH	Rser=39.5mohm	
Lpri2	4a	3	9.1uH	Rser=39.5mohm	
Laux1	2	1	11.42uH	Rser=116mohm	
Lsec1	6	10	37uH	Rser=90mohm	
Lsec2	7	9	37uH	Rser=180mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2       1					
.param Cprm1=54.95pf					
.param Cprm2=56.25pf					
.param Rdmp1=14505.8ohm					
.param Rdmp2=14505.8ohm					
Cpri1	5	4	{Cprm1}	Rser=10mohm	
Cpri2	4	3	{Cprm2}	Rser=10mohm	
Rdmp1	5	4	{Rdmp1}		
Rdmp2	4	3	{Rdmp2}		
Rg3	5	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg8	3	0	20meg		
Rg9	1	0	20meg		
Rg11	6	0	20meg		
Rg12	7	0	20meg		
Rg19	10	0	20meg		
Rg20	9	0	20meg		
.ends					

.subckt	750313082		5  4  3  2  1  6  9  7  10		
.param RxLkg=1453.1ohm					
.param Leakage=0.375uh					
Rlkg	5	5a	{RxLkg/2}		
L_Lkg	5	5a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	4	4a	{RxLkg/2}		
L_Lkg2	4	4a	{Leakage/2}	Rser=0.01mohm	
Lpri1	5a	4	9.063uH	Rser=41mohm	
Lpri2	4a	3	9.063uH	Rser=28mohm	
Laux1	2	1	11.42uH	Rser=123mohm	
Lsec1	6	9	1.827uH	Rser=8.4mohm	
Lsec2	7	10	1.827uH	Rser=8.4mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2       1					
.param Cprm1=9pf					
.param Cprm2=9pf					
.param Rdmp1=35843.03ohm					
.param Rdmp2=35843.03ohm					
Cpri1	5	4	{Cprm1}	Rser=10mohm	
Cpri2	4	3	{Cprm2}	Rser=10mohm	
Rdmp1	5	4	{Rdmp1}		
Rdmp2	4	3	{Rdmp2}		
Rg3	5	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg8	3	0	20meg		
Rg9	1	0	20meg		
Rg11	6	0	20meg		
Rg12	7	0	20meg		
Rg19	9	0	20meg		
Rg20	10	0	20meg		
.ends					

.subckt	750314433		2  5  1  3  4  10  7  6		
.param RxLkg=1748.02ohm					
.param Leakage=1.1uh					
Rlkg	2	2a	{RxLkg/2}		
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	5	5a	{RxLkg/2}		
L_Lkg2	5	5a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	5	44.45uH	Rser=154mohm	
Lpri2	5a	1	44.45uH	Rser=125mohm	
Laux1	3	4	23.472uH	Rser=230mohm	
Lsec1	10	7	5uH	Rser=10mohm	
Lsec2	7	6	5uH	Rser=148mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2       1					
.param Cprm1=11pf					
.param Cprm2=11pf					
.param Rdmp1=71509.75ohm					
.param Rdmp2=71509.75ohm					
Cpri1	2	5	{Cprm1}	Rser=10mohm	
Cpri2	5	1	{Cprm2}	Rser=10mohm	
Rdmp1	2	5	{Rdmp1}		
Rdmp2	5	1	{Rdmp2}		
Rg3	2	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg8	1	0	20meg		
Rg9	4	0	20meg		
Rg11	10	0	20meg		
Rg19	7	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt	750310035		3  4  2  1  7  9		
.param RxLkg=867.01ohm					
.param Leakage=0.8uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	76.6uH	Rser=87mohm	
Laux1	2	1	35.981uH	Rser=225mohm	
Lsec1	7	9	5.757uH	Rser=6mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=27.5pf					
.param Rdmp1=83883.14ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	7	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt	750032173		3  4  2  1  7  9		
.param RxLkg=6527.47ohm					
.param Leakage=6.75uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	120.25uH	Rser=480mohm	
Laux1	2	1	5.512uH	Rser=94mohm	
Lsec1	7	9	10.804uH	Rser=55mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=21.05pf					
.param Rdmp1=122813.13ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	7	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt	750310377		8  7  9  10  4  1		
.param RxLkg=469.69ohm					
.param Leakage=0.65uh					
Rlkg	8	8a	{RxLkg}		
L_Lkg	8	8a	{Leakage}	Rser=0.01mohm	
Lpri1	8a	7	126.35uH	Rser=180mohm	
Laux1	9	10	31.75uH	Rser=220mohm	
Lsec1	4	1	31.75uH	Rser=47.5mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=37.7pf					
.param Rdmp1=91769.91ohm					
Cpri1	8	7	{Cprm1}	Rser=10mohm	
Rdmp1	8	7	{Rdmp1}		
Rg3	8	0	20meg		
Rg5	9	0	20meg		
Rg7	7	0	20meg		
Rg9	10	0	20meg		
Rg11	4	0	20meg		
Rg19	1	0	20meg		
.ends					

.subckt	750310007		3  4  2  1  6  7  9  10		
.param RxLkg=945.19ohm					
.param Leakage=0.781uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	126.219uH	Rser=180mohm	
Laux1	2	1	40.781uH	Rser=250mohm	
Lsec1	6	7	3.528uH	Rser=13mohm	
Lsec2	9	10	40.781uH	Rser=105mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=13.44pf					
.param Rdmp1=153699.14ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	6	0	20meg		
Rg12	9	0	20meg		
Rg19	7	0	20meg		
Rg20	10	0	20meg		
.ends					

.subckt	750032395		3  1  4  5  10  9  8  6		
.param RxLkg=5138.3ohm					
.param Leakage=3.5uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	33.5uH	Rser=62mohm	
Laux1	4	5	10.152uH	Rser=425mohm	
Lsec1	10	9	0.336uH	Rser=19mohm	
Lsec2	8	6	1.342uH	Rser=6mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=31.35pf					
.param Rdmp1=54319.15ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	4	0	20meg		
Rg7	1	0	20meg		
Rg9	5	0	20meg		
Rg11	10	0	20meg		
Rg12	8	0	20meg		
Rg19	9	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt	750310310		3  1  4  5  10  9  8  6		
.param RxLkg=7618.9ohm					
.param Leakage=5uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	32uH	Rser=62mohm	
Laux1	4	5	10.152uH	Rser=425mohm	
Lsec1	10	9	1.342uH	Rser=6mohm	
Lsec2	8	6	1.342uH	Rser=55mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=29.1pf					
.param Rdmp1=56379.83ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	4	0	20meg		
Rg7	1	0	20meg		
Rg9	5	0	20meg		
Rg11	10	0	20meg		
Rg12	8	0	20meg		
Rg19	9	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt	750310027		3  4  2  1  5  7		
.param RxLkg=4681.68ohm					
.param Leakage=1.35uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	19.05uH	Rser=72mohm	
Laux1	2	1	6.296uH	Rser=135mohm	
Lsec1	5	7	1.007uH	Rser=6.75mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=10.19pf					
.param Rdmp1=70745.36ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	5	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310032		3  4  2  1  5  7		
.param RxLkg=2387.26ohm					
.param Leakage=4.5uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	150.5uH	Rser=390mohm	
Laux1	2	1	73.262uH	Rser=730mohm	
Lsec1	5	7	73.262uH	Rser=210mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=57.31pf					
.param Rdmp1=82227.79ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	5	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310031		3  4  2  1  5  7		
.param RxLkg=5138.95ohm					
.param Leakage=7.5uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	256.5uH	Rser=702mohm	
Laux1	2	1	10.995uH	Rser=50mohm	
Lsec1	5	7	21.551uH	Rser=40mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=20.17pf					
.param Rdmp1=180891.2ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	5	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310002		4  2  1  6  5  7  10		
.param RxLkg=655.38ohm					
.param Leakage=0.2uh					
Rlkg	4	4a	{RxLkg/2}		
L_Lkg	4	4a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}		
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	4a	2	6.9uH	Rser=13.5mohm	
Lpri2	2a	1	6.9uH	Rser=13.5mohm	
Laux1	6	5	17.286uH	Rser=105mohm	
Lsec1	7	10	2.286uH	Rser=8mohm	
K Lpri1 Lpri2 Laux1  Lsec1        1					
.param Cprm1=16.63pf					
.param Cprm2=16.4pf					
.param Rdmp1=22938.13ohm					
.param Rdmp2=22938.13ohm					
Cpri1	4	2	{Cprm1}	Rser=10mohm	
Cpri2	2	1	{Cprm2}	Rser=10mohm	
Rdmp1	4	2	{Rdmp1}		
Rdmp2	2	1	{Rdmp2}		
Rg3	4	0	20meg		
Rg5	6	0	20meg		
Rg7	2	0	20meg		
Rg8	1	0	20meg		
Rg9	5	0	20meg		
Rg11	7	0	20meg		
Rg19	10	0	20meg		
.ends					

.subckt	749119133		1  3  5  6  12  7  11  8  10  9		
.param RxLkg=2357.02ohm					
.param Leakage=2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	398uH	Rser=800mohm	
Laux1	5	6	25uH	Rser=600mohm	
Lsec1	12	7	2.778uH	Rser=20mohm	
Lsec2	11	8	2.778uH	Rser=20mohm	
Lsec3	10	9	2.778uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=4.5pf					
.param Rdmp1=471404.77ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg13	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
Rg21	9	0	20meg		
.ends					

.subckt	749119150		1  3  5  6  12  7  11  8  10  9		
.param RxLkg=2132.01ohm					
.param Leakage=2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	398uH	Rser=800mohm	
Laux1	5	6	25uH	Rser=500mohm	
Lsec1	12	7	7.716uH	Rser=60mohm	
Lsec2	11	8	7.716uH	Rser=60mohm	
Lsec3	10	9	7.716uH	Rser=60mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=5.5pf					
.param Rdmp1=426402.09ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg13	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
Rg21	9	0	20meg		
.ends					

.subckt	749119218		1  3  5  6  12  7  11  8  10  9		
.param RxLkg=5147.91ohm					
.param Leakage=3.2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	206.8uH	Rser=400mohm	
Laux1	5	6	23.333uH	Rser=800mohm	
Lsec1	12	7	0.771uH	Rser=7mohm	
Lsec2	11	8	0.771uH	Rser=7mohm	
Lsec3	10	9	0.771uH	Rser=7mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=4.6pf					
.param Rdmp1=337831.54ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg13	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
Rg21	9	0	20meg		
.ends					

.subckt	749119233		1  3  5  6  12  7  10  8		
.param RxLkg=3585.68ohm					
.param Leakage=1.8uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	208.2uH	Rser=200mohm	
Laux1	5	6	13.125uH	Rser=100mohm	
Lsec1	12	7	1.458uH	Rser=5mohm	
Lsec2	10	8	1.458uH	Rser=5mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=3pf					
.param Rdmp1=418329.7ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
.ends					

.subckt	749119250		1  3  5  6  12  7  11  8  10  9		
.param RxLkg=3161.68ohm					
.param Leakage=2.3uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	207.7uH	Rser=200mohm	
Laux1	5	6	17.865uH	Rser=100mohm	
Lsec1	12	7	5.833uH	Rser=30mohm	
Lsec2	11	8	5.833uH	Rser=30mohm	
Lsec3	10	9	5.833uH	Rser=30mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=6.3pf					
.param Rdmp1=288674.73ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg13	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
Rg21	9	0	20meg		
.ends					

.subckt	749119318		1  3  5  6  12  7  11  8  10  9		
.param RxLkg=2016.4ohm					
.param Leakage=1.1uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	118.9uH	Rser=100mohm	
Laux1	5	6	18.52uH	Rser=200mohm	
Lsec1	12	7	0.612uH	Rser=6mohm	
Lsec2	11	8	0.612uH	Rser=6mohm	
Lsec3	10	9	0.612uH	Rser=6mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=6.2pf					
.param Rdmp1=219970.55ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg13	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
Rg21	9	0	20meg		
.ends					

.subckt	749119333		1  3  5  6  12  7  11  8  10  9		
.param RxLkg=3194.49ohm					
.param Leakage=1.7uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	118.3uH	Rser=200mohm	
Laux1	5	6	7.5uH	Rser=100mohm	
Lsec1	12	7	0.833uH	Rser=10mohm	
Lsec2	11	8	0.833uH	Rser=10mohm	
Lsec3	10	9	0.833uH	Rser=10mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=5.9pf					
.param Rdmp1=225493.47ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg13	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
Rg21	9	0	20meg		
.ends					

.subckt	749119350		1  3  5  6  12  7  11  8  10  9		
.param RxLkg=2672.61ohm					
.param Leakage=1.2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	118.8uH	Rser=200mohm	
Laux1	5	6	7.5uH	Rser=100mohm	
Lsec1	12	7	2.315uH	Rser=20mohm	
Lsec2	11	8	2.315uH	Rser=20mohm	
Lsec3	10	9	2.315uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=4.2pf					
.param Rdmp1=267261.07ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg13	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
Rg21	9	0	20meg		
.ends					

.subckt	749119933		3  4  2  1  7  10  8  9		
.param RxLkg=692.1ohm					
.param Leakage=0.73uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	126.27uH	Rser=200mohm	
Laux1	2	1	31.75uH	Rser=300mohm	
Lsec1	7	10	3.528uH	Rser=20mohm	
Lsec2	8	9	3.528uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=21.9pf					
.param Rdmp1=120406.46ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg19	10	0	20meg		
Rg20	9	0	20meg
.ends					

.subckt	749119950		3  4  2  1  7  10  8  9		
.param RxLkg=2381.03ohm					
.param Leakage=1.2uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	125.8uH	Rser=200mohm	
Laux1	2	1	127uH	Rser=470mohm	
Lsec1	7	10	31.75uH	Rser=30mohm	
Lsec2	8	9	31.75uH	Rser=30mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=5pf					
.param Rdmp1=251992.41ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg19	10	0	20meg		
Rg20	9	0	20meg		
.ends					

.subckt	7491192912		1  3  5  6  12  10  8  7		
.param RxLkg=1606.04ohm					
.param Leakage=1.3uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	208.7uH	Rser=300mohm	
Laux1	5	6	36.458uH	Rser=200mohm	
Lsec1	12	10	3.281uH	Rser=20mohm	
Lsec2	10	8	1.458uH	Rser=10mohm	
Lsec3	8	7	17.865uH	Rser=60mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=7.8pf					
.param Rdmp1=259436.62ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg19	10	0	20meg		
Rg20	8	0	20meg		
Rg21	7	0	20meg		
.ends					

.subckt	7491193912		1  3  5  6  12  10  8  7		
.param RxLkg=1020.62ohm					
.param Leakage=0.5uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	119.5uH	Rser=200mohm	
Laux1	5	6	13.333uH	Rser=200mohm	
Lsec1	12	10	1.2uH	Rser=10mohm	
Lsec2	10	8	0.533uH	Rser=7mohm	
Lsec3	8	7	4.8uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=5pf					
.param Rdmp1=244949.23ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg19	10	0	20meg		
Rg20	8	0	20meg		
Rg21	7	0	20meg		
.ends					

.subckt	7491199112		3  4  2  1  7  10  8  9		
.param RxLkg=355.73ohm					
.param Leakage=0.3uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	126.7uH	Rser=200mohm	
Laux1	2	1	31.75uH	Rser=400mohm	
Lsec1	7	10	31.75uH	Rser=100mohm	
Lsec2	8	9	31.75uH	Rser=100mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=14pf					
.param Rdmp1=150594.26ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg19	10	0	20meg		
Rg20	9	0	20meg		
.ends					

.subckt	7491199212		3  4  2  1  7  10  8  9		
.param RxLkg=2312.66ohm					
.param Leakage=1.2uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	125.8uH	Rser=400mohm	
Laux1	2	1	31.75uH	Rser=90mohm	
Lsec1	7	10	31.75uH	Rser=40mohm	
Lsec2	8	9	31.75uH	Rser=40mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=5.3pf					
.param Rdmp1=244756.47ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg19	10	0	20meg		
Rg20	9	0	20meg		
.ends					

.subckt	7491199312		2  1  7  9		
.param RxLkg=294.63ohm					
.param Leakage=0.335uh					
Rlkg	2	2a	{RxLkg}		
L_Lkg	2	2a	{Leakage}	Rser=0.01mohm	
Lpri1	2a	1	39.665uH	Rser=99mohm	
Lsec1	7	9	40uH	Rser=63mohm	
K Lpri1    Lsec1        1					
.param Cprm1=80.8pf					
.param Rdmp1=35179.81ohm					
Cpri1	2	1	{Cprm1}	Rser=10mohm	
Rdmp1	2	1	{Rdmp1}		
Rg3	2	0	20meg		
Rg7	1	0	20meg		
Rg11	7	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt	7491199331		3  4  2  1  7  10  8  9		
.param RxLkg=3373.13ohm					
.param Leakage=1.7uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	125.3uH	Rser=400mohm	
Laux1	2	1	5.512uH	Rser=80mohm	
Lsec1	7	10	0.882uH	Rser=10mohm	
Lsec2	8	9	0.882uH	Rser=10mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=5pf					
.param Rdmp1=251992.41ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg19	10	0	20meg		
Rg20	9	0	20meg		
.ends					

.subckt	7491199332		1  2  5  4  7  8  9  6  10		
.param RxLkg=1318.37ohm					
.param Leakage=0.73uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	2	34.27uH	Rser=49mohm	
Laux1	5	4	8.75uH	Rser=180mohm	
Lsec1	7	8	0.432uH	Rser=69mohm	
Lsec2	8	9	0.972uH	Rser=11mohm	
Lsec3	6	10	2.701uH	Rser=14mohm	
K Lpri1  Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=21.9pf					
.param Rdmp1=63209.38ohm					
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	2	0	20meg		
Rg9	4	0	20meg		
Rg11	7	0	20meg		
Rg13	6	0	20meg		
Rg19	8	0	20meg		
Rg20	9	0	20meg		
Rg21	10	0	20meg		
.ends					

.subckt	7491199501		3  4  2  1  7  10  8  9		
.param RxLkg=2381.03ohm					
.param Leakage=1.2uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	125.8uH	Rser=400mohm	
Laux1	2	1	5.512uH	Rser=80mohm	
Lsec1	7	10	1.984uH	Rser=20mohm	
Lsec2	8	9	1.984uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=5pf					
.param Rdmp1=251992.41ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg9	1	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg19	10	0	20meg		
Rg20	9	0	20meg		
.ends					

.subckt	750310013		3  4  7  9		
.param RxLkg=513.38ohm					
.param Leakage=0.74uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	126.26uH	Rser=159mohm	
Lsec1	7	9	7.938uH	Rser=14mohm	
K Lpri1    Lsec1        1					
.param Cprm1=40.9pf					
.param Rdmp1=88107.25ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	7	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt	750310062		3  4  5  7		
.param RxLkg=1703.43ohm					
.param Leakage=2.5uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	4	124.5uH	Rser=456mohm	
Lsec1	5	7	7.938uH	Rser=22mohm	
K Lpri1    Lsec1        1					
.param Cprm1=42.4pf					
.param Rdmp1=86534.47ohm					
Cpri1	3	4	{Cprm1}	Rser=10mohm	
Rdmp1	3	4	{Rdmp1}		
Rg3	3	0	20meg		
Rg7	4	0	20meg		
Rg11	5	0	20meg		
Rg19	7	0	20meg		
.ends					


**********************************
************ WE-PoE+ **************
.subckt	750316333		1  3  4  5  8  6		
.param RxLkg=2269.9ohm					
.param Leakage=1.3uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	39.7uH	Rser=50mohm	
Laux1	4	5	5.766uH	Rser=89mohm	
Lsec1	8	6	5.766uH	Rser=13mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=20pf					
.param Rdmp1=71589.21ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt	750316332		1  3  4  5  8  6		
.param RxLkg=2886.75ohm					
.param Leakage=1.6uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	46.4uH	Rser=65mohm	
Laux1	4	5	9.293uH	Rser=140mohm	
Lsec1	8	6	1.92uH	Rser=5mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=16pf					
.param Rdmp1=86602.4ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt	750316331		1  3  4  5  8  6		
.param RxLkg=1326.83ohm					
.param Leakage=0.85uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	53.15uH	Rser=120mohm	
Laux1	4	5	11.344uH	Rser=125mohm	
Lsec1	8	6	0.844uH	Rser=4mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=19pf					
.param Rdmp1=84292.69ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt	750314783		5  4  3  2  1  6  9  7  10		
.param RxLkg=1736.83ohm					
.param Leakage=0.4uh					
Rlkg	5	5a	{RxLkg/2}		
L_Lkg	5	5a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	4	4a	{RxLkg/2}		
L_Lkg2	4	4a	{Leakage/2}	Rser=0.01mohm	
Lpri1	5a	4	6.3uH	Rser=47mohm	
Lpri2	4a	3	6.3uH	Rser=47mohm	
Laux1	2	1	8.025uH	Rser=233mohm	
Lsec1	6	9	1.284uH	Rser=8mohm	
Lsec2	7	10	1.284uH	Rser=8mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2       1					
.param Cprm1=10.2pf					
.param Cprm2=10.2pf					
.param Rdmp1=28223.54ohm					
.param Rdmp2=28223.54ohm					
Cpri1	5	4	{Cprm1}	Rser=10mohm	
Cpri2	4	3	{Cprm2}	Rser=10mohm	
Rdmp1	5	4	{Rdmp1}		
Rdmp2	4	3	{Rdmp2}		
Rg3	5	0	20meg		
Rg5	2	0	20meg		
Rg7	4	0	20meg		
Rg8	3	0	20meg		
Rg9	1	0	20meg		
Rg11	6	0	20meg		
Rg12	7	0	20meg		
Rg19	9	0	20meg		
Rg20	10	0	20meg		
.ends					

.subckt	750311320		1  2  4  5  6  9		
.param RxLkg=851.94ohm					
.param Leakage=0.6uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	2	99.4uH	Rser=100mohm	
Laux1	4	5	31.36uH	Rser=470mohm	
Lsec1	6	9	31.36uH	Rser=30mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=12.4pf					
.param Rdmp1=141990.56ohm					
Cpri1	1	2	{Cprm1}	Rser=10mohm	
Rdmp1	1	2	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	2	0	20meg		
Rg9	5	0	20meg		
Rg11	6	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt	750316116		1  3  5  6  11  7		
.param RxLkg=608.58ohm					
.param Leakage=0.2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	17.8uH	Rser=20mohm	
Laux1	5	6	4.5uH	Rser=66mohm	
Lsec1	11	7	4.5uH	Rser=11mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=15pf					
.param Rdmp1=54772.25ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	11	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310059		2  9  1  10  3  6		
.param RxLkg=8323.07ohm					
.param Leakage=1.5uh					
Rlkg	2	2a	{RxLkg}		
L_Lkg	2	2a	{Leakage}	Rser=0.01mohm	
Lpri1	2a	9	33.5uH	Rser=570mohm	
Laux1	1	10	6.699uH	Rser=530mohm	
Lsec1	3	6	0.547uH	Rser=2.8mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=2.32pf					
.param Rdmp1=194204.93ohm					
Cpri1	2	9	{Cprm1}	Rser=10mohm	
Rdmp1	2	9	{Rdmp1}		
Rg3	2	0	20meg		
Rg5	1	0	20meg		
Rg7	9	0	20meg		
Rg9	10	0	20meg		
Rg11	3	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt	750310167		1  3  2  4  5  6  12  11  10  9  8  7		
.param RxLkg=1440.05ohm					
.param Leakage=0.45uh					
Rlkg	1	1a	{RxLkg/2}		
L_Lkg	1	1a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg/2}		
L_Lkg2	2	2a	{Leakage/2}	Rser=0.01mohm	
Lpri1	1a	3	6.025uH	Rser=32mohm	
Lpri2	2a	4	6.025uH	Rser=32mohm	
Laux1	5	6	4uH	Rser=280mohm	
Lsec1	12	11	0.563uH	Rser=8.1mohm	
Lsec2	10	9	4uH	Rser=20.5mohm	
Lsec3	8	7	1uH	Rser=38mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=19.53pf					
.param Cprm2=21pf					
.param Rdmp1=20000.64ohm					
.param Rdmp2=20000.64ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Cpri2	2	4	{Cprm2}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rdmp2	2	4	{Rdmp2}		
Rg3	1	0	20meg		
Rg4	2	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg8	4	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	10	0	20meg		
Rg13	8	0	20meg		
Rg19	11	0	20meg		
Rg20	9	0	20meg		
Rg21	7	0	20meg		
.ends					

.subckt	750310346		1  3  2  4  5  6  12  7  11  8  10  9		
.param RxLkg=605.01ohm					
.param Leakage=1uh					
Rlkg	1	1a	{RxLkg*2}		
L_Lkg	1	1a	{Leakage*2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg*2}		
L_Lkg2	2	2a	{Leakage*2}	Rser=0.01mohm	
Lpri1	1a	3	99uH	Rser=221.2mohm	
Lpri2	2a	4	99uH	Rser=185.1mohm	
Laux1	5	6	11.111uH	Rser=245mohm	
Lsec1	12	7	11.111uH	Rser=66.4mohm	
Lsec2	11	8	11.111uH	Rser=68.9mohm	
Lsec3	10	9	11.111uH	Rser=68.7mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=34.15pf					
.param Cprm2=35.33pf					
.param Rdmp1=60500.79ohm					
.param Rdmp2=60500.79ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Cpri2	2	4	{Cprm2}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rdmp2	2	4	{Rdmp2}		
Rg3	1	0	20meg		
Rg4	2	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg8	4	0	20meg		
Rg9	6	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg13	10	0	20meg		
Rg19	7	0	20meg		
Rg20	8	0	20meg		
Rg21	9	0	20meg		
.ends					

.subckt	750310744		5  3  2  1  6  9		
.param RxLkg=2294.16ohm					
.param Leakage=0.6uh					
Rlkg	5	5a	{RxLkg}		
L_Lkg	5	5a	{Leakage}	Rser=0.01mohm	
Lpri1	5a	3	37.4uH	Rser=90mohm	
Laux1	2	1	38uH	Rser=200mohm	
Lsec1	6	9	6.08uH	Rser=3mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=4.5pf					
.param Rdmp1=145296.6ohm					
Cpri1	5	3	{Cprm1}	Rser=10mohm	
Rdmp1	5	3	{Rdmp1}		
Rg3	5	0	20meg		
Rg5	2	0	20meg		
Rg7	3	0	20meg		
Rg9	1	0	20meg		
Rg11	6	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt	750310743		5  3  2  1  6  9		
.param RxLkg=2019.71ohm					
.param Leakage=0.625uh					
Rlkg	5	5a	{RxLkg}		
L_Lkg	5	5a	{Leakage}	Rser=0.01mohm	
Lpri1	5a	3	37.375uH	Rser=82mohm	
Laux1	2	1	13.68uH	Rser=160mohm	
Lsec1	6	9	0.855uH	Rser=2mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=6.3pf					
.param Rdmp1=122798.15ohm					
Cpri1	5	3	{Cprm1}	Rser=10mohm	
Rdmp1	5	3	{Rdmp1}		
Rg3	5	0	20meg		
Rg5	2	0	20meg		
Rg7	3	0	20meg		
Rg9	1	0	20meg		
Rg11	6	0	20meg		
Rg19	9	0	20meg		
.ends					

.subckt	750310742		5  3  2  1  6  10		
.param RxLkg=1908.49ohm					
.param Leakage=0.47uh					
Rlkg	5	5a	{RxLkg}		
L_Lkg	5	5a	{Leakage}	Rser=0.01mohm	
Lpri1	5a	3	37.53uH	Rser=85mohm	
Laux1	2	1	11.495uH	Rser=155mohm	
Lsec1	6	10	9.5uH	Rser=25mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=3.99pf					
.param Rdmp1=154303.38ohm					
Cpri1	5	3	{Cprm1}	Rser=10mohm	
Rdmp1	5	3	{Rdmp1}		
Rg3	5	0	20meg		
Rg5	2	0	20meg		
Rg7	3	0	20meg		
Rg9	1	0	20meg		
Rg11	6	0	20meg		
Rg19	10	0	20meg		
.ends					

.subckt	750310927		3  1  5  6  7  8		
.param RxLkg=527.41ohm					
.param Leakage=0.9uh					
Rlkg	3	3a	{RxLkg}		
L_Lkg	3	3a	{Leakage}	Rser=0.01mohm	
Lpri1	3a	1	111.1uH	Rser=100mohm	
Laux1	5	6	3.111uH	Rser=60mohm	
Lsec1	7	8	12.444uH	Rser=50mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=65pf					
.param Rdmp1=65632.85ohm					
Cpri1	3	1	{Cprm1}	Rser=10mohm	
Rdmp1	3	1	{Rdmp1}		
Rg3	3	0	20meg		
Rg5	5	0	20meg		
Rg7	1	0	20meg		
Rg9	6	0	20meg		
Rg11	7	0	20meg		
Rg19	8	0	20meg		
.ends					

.subckt	7491194912		1  3  5  6  10  7		
.param RxLkg=515.95ohm					
.param Leakage=0.5uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	41.5uH	Rser=60mohm	
Laux1	5	6	4.667uH	Rser=180mohm	
Lsec1	10	7	4.667uH	Rser=18mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=55.9pf					
.param Rdmp1=43340.07ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	10	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310926		1  3  5  6  7  8  11  12		
.param RxLkg=570.54ohm					
.param Leakage=0.5uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	39.5uH	Rser=40mohm	
Laux1	5	6	2.5uH	Rser=200mohm	
Lsec1	7	8	1.6uH	Rser=9mohm	
Lsec2	11	12	2.5uH	Rser=200mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=48pf					
.param Rdmp1=45643.57ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	7	0	20meg		
Rg12	11	0	20meg		
Rg19	8	0	20meg		
Rg20	12	0	20meg		
.ends					

.subckt	749119450		1  3  5  6  10  7		
.param RxLkg=625.59ohm					
.param Leakage=0.8uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	64.3uH	Rser=100mohm	
Laux1	5	6	11.957uH	Rser=200mohm	
Lsec1	10	7	1.329uH	Rser=3mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=62.8pf					
.param Rdmp1=50907.31ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	10	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	7491194501		1  3  5  6  10  7		
.param RxLkg=765.56ohm					
.param Leakage=0.8uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	41.2uH	Rser=90mohm	
Laux1	5	6	4.339uH	Rser=170mohm	
Lsec1	10	7	0.857uH	Rser=5mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=65pf					
.param Rdmp1=40191.81ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	10	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	749119433		1  3  5  6  10  7		
.param RxLkg=3401.55ohm					
.param Leakage=3uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	39uH	Rser=99mohm	
Laux1	5	6	3.857uH	Rser=220mohm	
Lsec1	10	7	0.347uH	Rser=3.2mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=46.3pf					
.param Rdmp1=47621.74ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	10	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750310925		1  3  5  6  7  8  11  12		
.param RxLkg=1049.42ohm					
.param Leakage=1.2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	55.8uH	Rser=60mohm	
Laux1	5	6	3.563uH	Rser=350mohm	
Lsec1	7	8	0.891uH	Rser=8mohm	
Lsec2	11	12	3.563uH	Rser=350mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=57.35pf					
.param Rdmp1=49847.22ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	7	0	20meg		
Rg12	11	0	20meg		
Rg19	8	0	20meg		
Rg20	12	0	20meg		
.ends					


**********************************
************ WE-PoE++ **************
.subckt	750319035		1  5  3  4  11  7		
.param RxLkg=887.56ohm					
.param Leakage=0.55uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	5	15.45uH	Rser=25mohm	
Laux1	3	4	4uH	Rser=227mohm	
Lsec1	11	7	0.735uH	Rser=5mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=60pf					
.param Rdmp1=25819.87ohm					
Cpri1	1	5	{Cprm1}	Rser=10mohm	
Rdmp1	1	5	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg9	4	0	20meg		
Rg11	11	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750316335		1  3  4  5  8  6		
.param RxLkg=614.19ohm					
.param Leakage=0.325uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	49.675uH	Rser=26mohm	
Laux1	4	5	17.014uH	Rser=130mohm	
Lsec1	8	6	3.125uH	Rser=3mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=14pf					
.param Rdmp1=94491.25ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt	750343576		2  4  3  5  1  6  7  10  8  11		
.param RxLkg=225.73ohm					
.param Leakage=0.2uh					
Rlkg	2	2a	{RxLkg/2}		
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}		
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	4	24.9uH	Rser=5.1mohm	
Lpri2	3a	5	24.9uH	Rser=5.1mohm	
Laux1	1	6	25uH	Rser=95mohm	
Lsec1	7	10	25uH	Rser=7.1mohm	
Lsec2	8	11	25uH	Rser=7.1mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2       1					
.param Cprm1=39.25pf					
.param Cprm2=39.75pf					
.param Rdmp1=28216.69ohm					
.param Rdmp2=28216.69ohm					
Cpri1	2	4	{Cprm1}	Rser=10mohm	
Cpri2	3	5	{Cprm2}	Rser=10mohm	
Rdmp1	2	4	{Rdmp1}		
Rdmp2	3	5	{Rdmp2}		
Rg3	2	0	20meg		
Rg4	3	0	20meg		
Rg5	1	0	20meg		
Rg7	4	0	20meg		
Rg8	5	0	20meg		
Rg9	6	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg19	10	0	20meg		
Rg20	11	0	20meg		
.ends					

.subckt	750343164		2  4  3  5  1  6  7  10  8  11		
.param RxLkg=176.7ohm					
.param Leakage=0.43uh					
Rlkg	2	2a	{RxLkg/2}		
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}		
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	4	78.535uH	Rser=5.2mohm	
Lpri2	3a	5	78.535uH	Rser=4.8mohm	
Laux1	1	6	123.047uH	Rser=160mohm	
Lsec1	7	10	4.922uH	Rser=0.75mohm	
Lsec2	8	11	4.922uH	Rser=0.42mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2       1					
.param Cprm1=94pf					
.param Cprm2=94pf					
.param Rdmp1=32360.47ohm					
.param Rdmp2=32360.47ohm					
Cpri1	2	4	{Cprm1}	Rser=10mohm	
Cpri2	3	5	{Cprm2}	Rser=10mohm	
Rdmp1	2	4	{Rdmp1}		
Rdmp2	3	5	{Rdmp2}		
Rg3	2	0	20meg		
Rg4	3	0	20meg		
Rg5	1	0	20meg		
Rg7	4	0	20meg		
Rg8	5	0	20meg		
Rg9	6	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg19	10	0	20meg		
Rg20	11	0	20meg		
.ends					

.subckt	750318938		1  3  5  6  7  10		
.param RxLkg=155.58ohm					
.param Leakage=0.6uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	559.4uH	Rser=61mohm	
Laux1	5	6	236.6uH	Rser=372mohm	
Lsec1	7	10	35uH	Rser=4mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=66.4pf					
.param Rdmp1=145204.92ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg9	6	0	20meg		
Rg11	7	0	20meg		
Rg19	10	0	20meg		
.ends					

.subckt	750313355		1  3  2  4  5  6  7  10  8  11  9  12		
.param RxLkg=426.47ohm					
.param Leakage=0.479uh					
Rlkg	1	1a	{RxLkg*2}		
L_Lkg	1	1a	{Leakage*2}	Rser=0.01mohm	
Rlkg2	2	2a	{RxLkg*2}		
L_Lkg2	2	2a	{Leakage*2}	Rser=0.01mohm	
Lpri1	1a	3	99.521uH	Rser=102mohm	
Lpri2	2a	4	99.521uH	Rser=102mohm	
Laux1	5	6	25uH	Rser=229mohm	
Lsec1	7	10	25uH	Rser=33mohm	
Lsec2	8	11	25uH	Rser=33mohm	
Lsec3	9	12	25uH	Rser=33mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2 Lsec3      1					
.param Cprm1=15.7687pf					
.param Cprm2=15.7802pf					
.param Rdmp1=89033.99ohm					
.param Rdmp2=89033.99ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Cpri2	2	4	{Cprm2}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rdmp2	2	4	{Rdmp2}		
Rg3	1	0	20meg		
Rg4	2	0	20meg		
Rg5	5	0	20meg		
Rg7	3	0	20meg		
Rg8	4	0	20meg		
Rg9	6	0	20meg		
Rg11	7	0	20meg		
Rg12	8	0	20meg		
Rg13	9	0	20meg		
Rg19	10	0	20meg		
Rg20	11	0	20meg		
Rg21	12	0	20meg		
.ends					

.subckt	750310042		2  3  1  4  5  6  7  8		
.param RxLkg=1100.96ohm					
.param Leakage=2uh					
Rlkg	2	2a	{RxLkg}		
L_Lkg	2	2a	{Leakage}	Rser=0.01mohm	
Lpri1	2a	3	273uH	Rser=40mohm	
Laux1	1	4	68.75uH	Rser=50mohm	
Lsec1	5	6	68.75uH	Rser=10mohm	
Lsec2	7	8	68.75uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=30pf					
.param Rdmp1=151382.67ohm					
Cpri1	2	3	{Cprm1}	Rser=10mohm	
Rdmp1	2	3	{Rdmp1}		
Rg3	2	0	20meg		
Rg5	1	0	20meg		
Rg7	3	0	20meg		
Rg9	4	0	20meg		
Rg11	5	0	20meg		
Rg12	7	0	20meg		
Rg19	6	0	20meg		
Rg20	8	0	20meg		
.ends					

.subckt	750316336		1  3  4  5  8  6		
.param RxLkg=651.77ohm					
.param Leakage=0.47uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	49.53uH	Rser=14mohm	
Laux1	4	5	12.5uH	Rser=62mohm	
Lsec1	8	6	12.5uH	Rser=8mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=26pf					
.param Rdmp1=69337.46ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt	750316334		1  3  4  5  8  6		
.param RxLkg=816.67ohm					
.param Leakage=0.49uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	49.51uH	Rser=25mohm	
Laux1	4	5	12.5uH	Rser=83mohm	
Lsec1	8	6	1.02uH	Rser=3mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=18pf					
.param Rdmp1=83333.26ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	8	0	20meg		
Rg19	6	0	20meg		
.ends					

.subckt	750313095		2  4  3  5  1  6  8  12  7  11		
.param RxLkg=566.06ohm					
.param Leakage=0.5uh					
Rlkg	2	2a	{RxLkg/2}		
L_Lkg	2	2a	{Leakage/2}	Rser=0.01mohm	
Rlkg2	3	3a	{RxLkg/2}		
L_Lkg2	3	3a	{Leakage/2}	Rser=0.01mohm	
Lpri1	2a	4	61.475uH	Rser=19mohm	
Lpri2	3a	5	61.475uH	Rser=21.6mohm	
Laux1	1	6	102.035uH	Rser=188mohm	
Lsec1	8	12	20.155uH	Rser=13mohm	
Lsec2	7	11	20.155uH	Rser=12.6mohm	
K Lpri1 Lpri2 Laux1  Lsec1 Lsec2       1					
.param Cprm1=15.8pf					
.param Cprm2=15.8pf					
.param Rdmp1=69880.69ohm					
.param Rdmp2=69880.69ohm					
Cpri1	2	4	{Cprm1}	Rser=10mohm	
Cpri2	3	5	{Cprm2}	Rser=10mohm	
Rdmp1	2	4	{Rdmp1}		
Rdmp2	3	5	{Rdmp2}		
Rg3	2	0	20meg		
Rg4	3	0	20meg		
Rg5	1	0	20meg		
Rg7	4	0	20meg		
Rg8	5	0	20meg		
Rg9	6	0	20meg		
Rg11	8	0	20meg		
Rg12	7	0	20meg		
Rg19	12	0	20meg		
Rg20	11	0	20meg		
.ends					

.subckt	750318961		1  5  3  4  11  7		
.param RxLkg=161.37ohm					
.param Leakage=0.25uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	5	99.75uH	Rser=12.7mohm	
Laux1	3	4	39.063uH	Rser=80mohm	
Lsec1	11	7	6.25uH	Rser=2mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=60pf					
.param Rdmp1=64549.68ohm					
Cpri1	1	5	{Cprm1}	Rser=10mohm	
Rdmp1	1	5	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg9	4	0	20meg		
Rg11	11	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750318962		1  5  3  4  12  9  10  7		
.param RxLkg=81.65ohm					
.param Leakage=0.2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	5	99.8uH	Rser=9mohm	
Laux1	3	4	39.063uH	Rser=68mohm	
Lsec1	12	9	39.063uH	Rser=10mohm	
Lsec2	10	7	39.063uH	Rser=10mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=150pf					
.param Rdmp1=40825ohm					
Cpri1	1	5	{Cprm1}	Rser=10mohm	
Rdmp1	1	5	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg9	4	0	20meg		
Rg11	12	0	20meg		
Rg12	10	0	20meg		
Rg19	9	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	750319020		1  5  3  4  11  7		
.param RxLkg=442.81ohm					
.param Leakage=0.4uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	5	16.6uH	Rser=11mohm	
Laux1	3	4	4.25uH	Rser=122mohm	
Lsec1	11	7	0.68uH	Rser=2mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=120pf					
.param Rdmp1=18819.26ohm					
Cpri1	1	5	{Cprm1}	Rser=10mohm	
Rdmp1	1	5	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg9	4	0	20meg		
Rg11	11	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750319021		1  5  3  4  10  7		
.param RxLkg=486.56ohm					
.param Leakage=0.5uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	5	21.5uH	Rser=12mohm	
Laux1	3	4	3.819uH	Rser=125mohm	
Lsec1	10	7	3.819uH	Rser=4mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=120pf					
.param Rdmp1=21408.66ohm					
Cpri1	1	5	{Cprm1}	Rser=10mohm	
Rdmp1	1	5	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg9	4	0	20meg		
Rg11	10	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750319032		1  5  3  4  11  7		
.param RxLkg=381.39ohm					
.param Leakage=0.48uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	5	21.52uH	Rser=12mohm	
Laux1	3	4	3.819uH	Rser=125mohm	
Lsec1	11	7	15.278uH	Rser=12mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=180pf					
.param Rdmp1=17480.16ohm					
Cpri1	1	5	{Cprm1}	Rser=10mohm	
Rdmp1	1	5	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg9	4	0	20meg		
Rg11	11	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750319033		1  6  3  4  10  7		
.param RxLkg=260.64ohm					
.param Leakage=0.25uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	6	99.75uH	Rser=11mohm	
Laux1	3	4	39.063uH	Rser=51mohm	
Lsec1	10	7	6.25uH	Rser=2mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=23pf					
.param Rdmp1=104256.89ohm					
Cpri1	1	6	{Cprm1}	Rser=10mohm	
Rdmp1	1	6	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	6	0	20meg		
Rg9	4	0	20meg		
Rg11	10	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750319034		1  6  3  4  12  9  11  8		
.param RxLkg=73.03ohm					
.param Leakage=0.16uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	6	99.84uH	Rser=11mohm	
Laux1	3	4	39.063uH	Rser=51mohm	
Lsec1	12	9	39.063uH	Rser=9mohm	
Lsec2	11	8	39.063uH	Rser=9mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=120pf					
.param Rdmp1=45643.57ohm					
Cpri1	1	6	{Cprm1}	Rser=10mohm	
Rdmp1	1	6	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	6	0	20meg		
Rg9	4	0	20meg		
Rg11	12	0	20meg		
Rg12	11	0	20meg		
Rg19	9	0	20meg		
Rg20	8	0	20meg		
.ends					

.subckt	750319036		1  5  3  4  10  7		
.param RxLkg=595.91ohm					
.param Leakage=0.5uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	5	15.5uH	Rser=24mohm	
Laux1	3	4	2.939uH	Rser=200mohm	
Lsec1	10	7	2.939uH	Rser=5mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=110pf					
.param Rdmp1=19069.22ohm					
Cpri1	1	5	{Cprm1}	Rser=10mohm	
Rdmp1	1	5	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg9	4	0	20meg		
Rg11	10	0	20meg		
Rg19	7	0	20meg		
.ends					

.subckt	750319069		1  5  3  4  11  7		
.param RxLkg=405.17ohm					
.param Leakage=0.41uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	5	15.59uH	Rser=22mohm	
Laux1	3	4	4uH	Rser=150mohm	
Lsec1	11	7	13.796uH	Rser=22mohm	
K Lpri1  Laux1  Lsec1        1					
.param Cprm1=160pf					
.param Rdmp1=15811.41ohm					
Cpri1	1	5	{Cprm1}	Rser=10mohm	
Rdmp1	1	5	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	3	0	20meg		
Rg7	5	0	20meg		
Rg9	4	0	20meg		
Rg11	11	0	20meg		
Rg19	7	0	20meg		
.ends					


**********************************
************ WE-PoEH **************
.subckt	749119550		1  3  4  5  9  6  10  7		
.param RxLkg=1242.26ohm					
.param Leakage=0.4uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	47.6uH	Rser=50mohm	
Laux1	4	5	6.75uH	Rser=80mohm	
Lsec1	9	6	1.688uH	Rser=7mohm	
Lsec2	10	7	1.688uH	Rser=7mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=5.4pf					
.param Rdmp1=149071.34ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491195331		1  3  4  5  9  6  10  7		
.param RxLkg=791.56ohm					
.param Leakage=0.2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	20.8uH	Rser=20mohm	
Laux1	4	5	11.813uH	Rser=120mohm	
Lsec1	9	6	1.313uH	Rser=7mohm	
Lsec2	10	7	1.313uH	Rser=7mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=7.6pf					
.param Rdmp1=83113.74ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	749119533		1  3  4  5  9  6  10  7		
.param RxLkg=1506.46ohm					
.param Leakage=0.5uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	53.5uH	Rser=50mohm	
Laux1	4	5	7.594uH	Rser=80mohm	
Lsec1	9	6	0.844uH	Rser=4mohm	
Lsec2	10	7	0.844uH	Rser=4mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=5.1pf					
.param Rdmp1=162697.98ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491195224		1  3  4  5  9  6  10  7		
.param RxLkg=344.06ohm					
.param Leakage=0.23uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	20.77uH	Rser=20mohm	
Laux1	4	5	9.333uH	Rser=110mohm	
Lsec1	9	6	47.25uH	Rser=110mohm	
Lsec2	10	7	47.25uH	Rser=110mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=53.2pf					
.param Rdmp1=31414.05ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491195212		1  3  4  5  9  6  10  7		
.param RxLkg=377.96ohm					
.param Leakage=0.12uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	20.88uH	Rser=25mohm	
Laux1	4	5	9.333uH	Rser=110mohm	
Lsec1	9	6	11.813uH	Rser=47mohm	
Lsec2	10	7	11.813uH	Rser=47mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=12pf					
.param Rdmp1=66143.79ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491195112		1  3  4  5  9  6  10  7		
.param RxLkg=879.16ohm					
.param Leakage=0.3uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	40.7uH	Rser=53mohm	
Laux1	4	5	5.766uH	Rser=83mohm	
Lsec1	9	6	5.766uH	Rser=16mohm	
Lsec2	10	7	5.766uH	Rser=19mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=7.1pf					
.param Rdmp1=120152.42ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491195501		1  3  4  5  9  6  10  7		
.param RxLkg=843.05ohm					
.param Leakage=0.2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	20.8uH	Rser=30mohm	
Laux1	4	5	9.333uH	Rser=110mohm	
Lsec1	9	6	2.333uH	Rser=10mohm	
Lsec2	10	7	2.333uH	Rser=10mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=6.7pf					
.param Rdmp1=88520.13ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491196212		1  3  4  5  9  6  10  7		
.param RxLkg=8.04ohm					
.param Leakage=0.02uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	127.98uH	Rser=10mohm	
Laux1	4	5	392uH	Rser=300mohm	
Lsec1	9	6	578uH	Rser=80mohm	
Lsec2	10	7	578uH	Rser=100mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=121pf					
.param Rdmp1=51426.01ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491196112		1  3  4  5  9  6  10  7		
.param RxLkg=307.15ohm					
.param Leakage=0.2uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	99.8uH	Rser=40mohm	
Laux1	4	5	25uH	Rser=80mohm	
Lsec1	9	6	34.028uH	Rser=20mohm	
Lsec2	10	7	34.028uH	Rser=30mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=10.6pf					
.param Rdmp1=153573.62ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491196501		1  3  4  5  9  6  10  7		
.param RxLkg=65.59ohm					
.param Leakage=0.1uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	127.9uH	Rser=10mohm	
Laux1	4	5	392uH	Rser=300mohm	
Lsec1	9	6	98uH	Rser=20mohm	
Lsec2	10	7	98uH	Rser=30mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=45.4pf					
.param Rdmp1=83955.42ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	749119650		1  3  4  5  9  6  10  7		
.param RxLkg=168.55ohm					
.param Leakage=0.1uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	99.9uH	Rser=30mohm	
Laux1	4	5	25uH	Rser=90mohm	
Lsec1	9	6	6.25uH	Rser=7mohm	
Lsec2	10	7	6.25uH	Rser=7mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=8.8pf					
.param Rdmp1=168550.22ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	7491196331		1  3  4  5  9  6  10  7		
.param RxLkg=454.75ohm					
.param Leakage=0.3uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	127.7uH	Rser=50mohm	
Laux1	4	5	98uH	Rser=300mohm	
Lsec1	9	6	12.5uH	Rser=10mohm	
Lsec2	10	7	12.5uH	Rser=10mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=8.5pf					
.param Rdmp1=194028.78ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt	749119633		1  3  4  5  9  6  10  7		
.param RxLkg=617.54ohm					
.param Leakage=0.3uh					
Rlkg	1	1a	{RxLkg}		
L_Lkg	1	1a	{Leakage}	Rser=0.01mohm	
Lpri1	1a	3	99.7uH	Rser=20mohm	
Laux1	4	5	25uH	Rser=80mohm	
Lsec1	9	6	2.778uH	Rser=6mohm	
Lsec2	10	7	2.778uH	Rser=6mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=5.9pf					
.param Rdmp1=205846.58ohm					
Cpri1	1	3	{Cprm1}	Rser=10mohm	
Rdmp1	1	3	{Rdmp1}		
Rg3	1	0	20meg		
Rg5	4	0	20meg		
Rg7	3	0	20meg		
Rg9	5	0	20meg		
Rg11	9	0	20meg		
Rg12	10	0	20meg		
Rg19	6	0	20meg		
Rg20	7	0	20meg		
.ends					
