**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Common Mode Power Line Choke
* Matchcode:              WE-CMB 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-26
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.SUBCKT CMB    1  2  3  4  PARAMS: 
R_R9  N12325  3  {R2}
R_R8  N13265  N13287  {Rs4}
Kn_K6  L_L11  L_L12  
+  L_L13  L_L14  0.9999
R_R3  N12571  N12583  {Rs3}
R_R10  N13777  4  {R2}
C_C10  N13029  N12821  {ck}
R_R20  N13215  N13229  {dR4}
L_L11  N12821  N12295  {dL4}
R_R17  N12267  N12273  {dR3}
L_L8  N13265  N13287  {L4}
R_R7  N13287  N13305  {Rs3}
L_L9  N12295  N12307  {L5}
Kn_K4  L_L7  L_L8  1
R_R2  N12583  N12599  {Rs2}
Kn_K5  L_L9  L_L10  1
R_R16  N13229  N13249  {dR6}
Kn_K7  L_L15  L_L16  
+  L_L17  L_L18  0.9999
C_C5  N12273  N12289  {dC4}
L_L6  N13287  N13305  {L3}
L_L7  N12307  N12571  {L4}
R_R6  N13305  N13319  {Rs2}
R_R21  1  N12257  {Rdc}
Kn_K3  L_L5  L_L6  1
L_L16  N12257  N12799  {dL3}
C_C8  N13215  N13741  {dC3}
L_L18  N13023  N13215  {dL3}
R_R1  N12599  3  {Rs1}
R_R13  N12289  N12295  {dR5}
L_L4  N13305  N13319  {L2}
L_L5  N12571  N12583  {L3}
R_R15  N13755  N13249  {dR5}
R_R5  N13319  4  {Rs1}
R_R18  N12257  N12273  {dR4}
Kn_K2  L_L3  L_L4  1
R_R19  N13741  N13229  {dR3}
L_L15  N12799  N12273  {dL3}
L_L17  N13229  N13023  {dL3}
L_L3  N12583  N12599  {L2}
R_R11  N12295  N12307  {Rs5}
L_L2  N13319  4  {L1}
C_C4  N13249  N13265  {C2}
L_L10  N13249  N13265  {L5}
Kn_K1  L_L1  L_L2  1
R_R14  N12273  N12295  {dR6}
C_C6  N13229  N13755  {dC4}
L_L12  N12273  N12821  {dL4}
L_L14  N13029  N13229  {dL4}
L_L1  N12599  3  {L1}
C_C1  N12307  N12325  {C1}
R_R12  N13249  N13265  {Rs5}
C_C2  N13265  N13777  {C1}
R_R22  2  N13215  {Rdc}
C_C9  N13023  N12799  {ck}
R_R4  N12307  N12571  {Rs4}
C_C3  N12295  N12307  {C2}
L_L13  N13249  N13029  {dL4}
C_C7  N12257  N12267  {dC3} 
.ends  CMB
****
.subckt CMB1 1 2 3 4 PARAMS:
+ L3=1150u
+ Rs3=6.4k
+ C1=12p
+ R2=1
+ L1=0.1p
+ Rs2=700
+ C2=0.1u
+ Rs1=10
+ L2=1u
+ L4=0.01u
+ Rs4=1
+ L5=0.01p
+ Rs5=0.1k
+ dR5=1
+ Rdc=1m
+ ck=3p
+ dR3=1k
+ dR6=2.8k
+ dR4=1k
+ dC3=2.1p
+ dL3=0.2u
+ dC4=1p
+ dL4=0.245u
L5 N009 N008 {L3}
C3 N002 N001 {C1}
L1 4 N010 {L1}
L3 N010 N009 {L2}
L6 N015 N014 {L3}
C4 N024 N013 {C1}
L2 3 N016 {L1}
L4 N016 N015 {L2}
L8 N014 N013 {L4}
L7 N008 N001 {L4}
L9 N001 N007 {L5}
L10 N013 N021 {L5}
R1 N003 1 {Rdc}
R2 N005 N003 {dR4}
C1 N004 N003 {dC3}
L17 N011 N003 {dL3}
L18 N017 N018 {dL3}
C2 N011 N018 {ck}
R3 N005 N004 {dR3}
R4 N019 N022 {dR3}
C9 N022 N017 {dC3}
R5 N019 N017 {dR4}
L19 N005 N011 {dL3}
L20 N018 N019 {dL3}
R6 N017 2 {Rdc}
R8 N007 N005 {dR6}
C10 N006 N005 {dC4}
L13 N012 N005 {dL4}
L14 N019 N020 {dL4}
C11 N012 N020 {ck}
R9 N007 N006 {dR5}
R10 N021 N023 {dR5}
C12 N023 N019 {dC4}
R11 N021 N019 {dR6}
L15 N007 N012 {dL4}
L16 N020 N021 {dL4}
R7 N001 N007 {Rs5}
C5 N001 N007 {C2}
R12 N013 N021 {Rs5}
C6 N013 N021 {C2}
R13 N008 N001 {Rs4}
R14 N009 N008 {Rs3}
R15 N010 N009 {Rs2}
R16 4 N010 {Rs1}
R17 N014 N013 {Rs4}
R18 N015 N014 {Rs3}
R19 N016 N015 {Rs2}
R20 3 N016 {Rs1}
R21 4 N002 {R2}
R22 3 N024 {R2}
K3 L5 L6 1
K2 L3 L4 1
K1 L1 L2 1
K4 L7 L8 1
K5 L9  L10 1
K7 L17 L18 L19 L20 0.9999
K6 L13 L14 L15 L16 0.9999
.ends
****
.subckt XS_744821201_1m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=7u
+  DL4=18n
+  DC3=0.2p 
+  DC4=10p 
+  DR3=7000
+  DR4=7000
+  DR5=60000
+  DR6=7000
+  Rdc=0.33
+  ck=40pF
+  L1=15m
+  L2=10u
+  L3=2n
+  L4=35n
+  L5=0.25n
+  C1=25p
+  C2=25p
+  RS1=200000
+  RS2=7000
+  RS3=5000
+  RS4=5000
+  RS5=4000
+  R2=0.08
.ends XS_744821201_1m
****
.subckt XS_744821240_4m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000017
+  DL4=0.000000035
+  DC3=0.000000000006
+  DC4=0.000000000003
+  DR3=17
+  dR4=11.25k
+  DR5=230
+  dR6=50k
+  Rdc=0.082
+  ck=2pF
+  L1=3.3m
+  L2=0.81m
+  L3=23u
+  L4=40u
+  L5=570.4n
+  C1=12.2p
+  C2=1
+  Rs1=19.5k
+  Rs2=29k
+  RS3=500
+  RS4=600
+  RS5=2000
+  R2=10.41
.ends XS_744821240_4m
****
.subckt XS_744821150_5m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000018
+  DL4=0.000000064
+  DC3=0.0000000000125
+  DC4=0.000000000005
+  DR3=17
+  dR4=15k
+  DR5=30
+  dR6=2k
+  Rdc=0.168
+  ck=2pF
+  L1=3.6m
+  L2=0.8m
+  L3=23u
+  L4=4u
+  L5=800.4n
+  C1=11.5p
+  C2=4p
+  Rs1=19k
+  Rs2=19k
+  RS3=500
+  RS4=200
+  RS5=2500
+  R2=1
.ends XS_744821150_5m
****
.subckt XS_744821110_10m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000052
+  DL4=0.000000005
+  DC3=0.000000000022
+  DC4=0.000000000006
+  DR3=17
+  dR4=25k
+  dR5=30k
+  dR6=5k
+  Rdc=0.266
+  ck=6pF
+  L1=8.8m
+  L2=0.180m
+  L3=23u
+  L4=4u
+  L5=520.4n
+  C1=14p
+  C2=10p
+  Rs1=69k
+  Rs2=20k
+  RS3=500
+  RS4=200
+  RS5=800
+  R2=1
.ends XS_744821110_10m
****
.subckt XS_744821120_20m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.000011
+  DL4=0.000000007
+  DC3=0.000000000019
+  DC4=0.000000000001
+  DR3=17
+  dR4=30k
+  DR5=30
+  dR6=8k
+  Rdc=0.779
+  ck=12pF
+  L1=19.8m
+  L2=1.8m
+  L3=23u
+  L4=4u
+  L5=2.920u
+  C1=11p
+  C2=15p
+  Rs1=129k
+  Rs2=20k
+  RS3=500
+  RS4=200
+  RS5=2200
+  R2=20.41
.ends XS_744821120_20m
****
.subckt XS_744821039_39m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.000022
+  DL4=0.000000225
+  DC3=0.000000000027
+  DC4=0.000000000038
+  DR3=17
+  dR4=127k
+  DR5=23
+  dR6=1.5k
+  Rdc=1.905
+  ck=3pF
+  L1=37.5m
+  L2=1.8m
+  L3=23u
+  L4=4u
+  L5=630n
+  C1=27p
+  C2=90p
+  Rs1=499k
+  Rs2=29k
+  RS3=500
+  RS4=200
+  RS5=1000
+  R2=1
.ends XS_744821039_39m
****
.subckt S_744822301_1m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=0.00060538
+  L2=0.00010035
+  L3=0.00004247
+  L4=0.00001022
+  L5=0.000000036
+  C1=0.000000000003
+  C2=0.000000000001
+  RS1=8828
+  RS2=1447
+  RS3=703
+  RS4=678
+  RS5=509
+  R2=0.11
+  DL3=0.00000031037
+  DL4=0.00000001106
+  DC3=0.00000000000019056
+  DC4=0.000000000007
+  DR3=1000
+  DR4=4500
+  DR5=11000
+  DR6=438
+  Rdc=0.021
+  ck=12.5pF
.ends S_744822301_1m
****
.subckt S_744822233_3.3m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000014
+  DL4=0.000000003
+  DC3=0.0000000000083
+  DC4=0.000000000002
+  DR3=17
+  dR4=22k
+  DR5=30
+  dR6=2k
+  Rdc=0.079
+  ck=3pF
+  L1=3m
+  L2=0.58m
+  L3=23u
+  L4=4u
+  L5=210.4n
+  C1=8p
+  C2=8p
+  Rs1=38k
+  Rs2=6k
+  RS3=500
+  RS4=200
+  RS5=1200
+  R2=1.41
.ends S_744822233_3.3m
****
.subckt S_744822110_10m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000035
+  DL4=0.000000104
+  DC3=0.0000000000192
+  DC4=0.000000000019
+  DR3=17
+  dR4=27k
+  DR5=30
+  dR6=12k
+  Rdc=0.236
+  ck=4pF
+  L1=11.6m
+  L2=800u
+  L3=23u
+  L4=4u
+  L5=1.8u
+  C1=14.5p
+  C2=8p
+  Rs1=79k
+  Rs2=19k
+  RS3=500
+  RS4=200
+  RS5=5000
+  R2=10.41
.ends S_744822110_10m
****
.subckt S_744822120_20m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000068
+  DL4=0.00000001
+  DC3=0.000000000032
+  DC4=0.000000000003
+  DR3=17
+  dR4=27k
+  DR5=30
+  dR6=2k
+  Rdc=0.355
+  ck=10pF
+  L1=16.6m
+  L2=800u
+  L3=23u
+  L4=4u
+  L5=80.4n
+  C1=26.5p
+  C2=28p
+  Rs1=340k
+  Rs2=19k
+  RS3=500
+  RS4=200
+  RS5=800
+  R2=1.41
.ends S_744822120_20m
****
.subckt M_744823305_5m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=0.0000149932488790583
+  L2=0.0000219946000050973
+  L3=0.0000734873979778146
+  L4=0.00545630375790193
+  L5=9.38962438216997E-10
+  C1=1.50319062754058E-11
+  C2=5.341200990649E-12
+  RS1=5265.31166846459
+  RS2=7902.70514846992
+  RS3=1651.19231206434
+  RS4=39361.136544689
+  RS5=9214.69726890499
+  R2=0.109490257696781
+  DL3=0.0000017
+  DL4=0.00000002
+  DC3=0.000000000033
+  DC4=0.00000000006
+  DR3=4
+  DR4=1120
+  DR5=6
+  DR6=800
+  Rdc=60.229m
+  ck=4pF
.ends M_744823305_5m
****
.subckt M_744823601_1m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.00000024233
+  DC3=0.00000000001
+  DL4=0.00000001079
+  DC4=0.00000000000421
+  DR3=10
+  DR4=3300
+  DR5=173
+  DR6=2705
+  Rdc=8.952m
+  ck=2.005pF
+  L1=0.00001849
+  L2=0.000039
+  L3=0.000019
+  L4=0.0009
+  L5=0.00000001869
+  C1=0.00000000000305
+  C2=0.00000000000415
+  RS1=745
+  RS2=200
+  RS3=332
+  RS4=3200
+  RS5=362
+  R2=11
.ends M_744823601_1m
****
.subckt M_744823422_2.2m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=3m
+  L2=800.72u
+  L3=523.19u
+  L4=242.84u
+  L5=42.11n
+  C1=3.43p
+  C2=4.39p
+  RS1=7554
+  RS2=1544
+  RS3=1544
+  RS4=2457
+  RS5=561
+  R2=39
+  dL3=532.17n
+  dC3=11.33p
+  dL4=27.79n
+  dC4=4.13p
+  DR3=28
+  DR4=10212
+  DR5=23
+  DR6=2190
+  Rdc=24.288m
+  ck=2p
.ends M_744823422_2.2m
****
.subckt M_744823333_3.3m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000008388
+  DC3=0.0000000000124
+  DL4=0.00000004038
+  DC4=0.00000000000673
+  DR3=0.21
+  DR4=7180
+  DR5=45
+  DR6=1197
+  Rdc=45.566m
+  ck=2.005pF
+  L1=2m
+  L2=0.00038766
+  L3=0.00021925
+  L4=0.007228
+  L5=0.000000082
+  C1=0.00000000000368
+  C2=0.00000000000359
+  RS1=549
+  RS2=539
+  RS3=539
+  RS4=18717
+  RS5=756
+  R2=39
.ends M_744823333_3.3m
****
.subckt M_744823210_10m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.00000268
+  DC3=0.000000000026
+  DL4=0.00000007674
+  DC4=0.000000000032
+  DR3=1.43
+  DR4=11000
+  DR5=0.019
+  DR6=1052
+  Rdc=99.542m
+  ck=2.005pF
+  L1=10m
+  L2=2m
+  L3=203u
+  L4=104u
+  L5=900.4n
+  C1=16.7p
+  C2=20p
+  Rs1=48k
+  Rs2=29k
+  Rs3=5k
+  Rs4=5k
+  Rs5=2k
+  R2=40.41
.ends M_744823210_10m
****
.subckt M_744823220_20m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000062
+  DL4=0.000000095
+  DC3=0.000000000032
+  DC4=0.00000000006
+  DR3=17
+  dR4=30k
+  DR5=23
+  dR6=4k
+  Rdc=216.759m
+  ck=3pF
+  L1=19m
+  L2=0.000059
+  L3=0.000092
+  L4=0.000021
+  L5=0.000000124
+  C1=0.000000000022
+  C2=0.00000000003
+  Rs1=124k
+  Rs2=199k
+  RS3=561
+  RS4=915
+  RS5=894
+  R2=1
.ends M_744823220_20m
****
.subckt L_744824101_1m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.00000040534
+  DC3=0.00000000001907
+  DL4=0.00000001675
+  DC4=0.00000000000382
+  DR3=10
+  DR4=4300
+  DR5=0.63
+  DR6=1750
+  Rdc=6.372m
+  ck=2.005pF
+  L1=0.00172384
+  L2=0.00089876
+  L3=0.00015148
+  L4=0.0001977
+  L5=0.0000001268
+  C1=0.00000000000832
+  C2=0.00000000000548
+  RS1=565
+  RS2=470
+  RS3=557
+  RS4=2992
+  RS5=643
+  R2=0.56
.ends L_744824101_1m
****
.subckt L_744824622_2.2m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.00000068242
+  DC3=0.00000000001367
+  DL4=0.000000029
+  DC4=0.00000000000971
+  DR3=0.02
+  DR4=6278
+  DR5=28
+  DR6=821
+  Rdc=16.345m
+  ck=2pF
+  L1=0.00000897
+  L2=0.00016374
+  L3=0.00013744
+  L4=0.00443191
+  L5=0.00000010639
+  C1=0.00000000000399
+  C2=0.00000000000211
+  RS1=10
+  RS2=943
+  RS3=928
+  RS4=8391
+  RS5=765
+  R2=4
.ends L_744824622_2.2m
****
.subckt L_744824433_3.3m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  dL3=1u
+  dL4=50.25n
+  dC3=15.595p
+  dC4=8.4p
+  DR3=0.1
+  dR4=8k
+  DR5=0.1
+  DR6=900
+  Rdc=28.429m
+  ck=2pF
+  L1=0.000001023
+  L2=0.00013929
+  L3=0.00017837
+  L4=0.00099218
+  L5=0.0000000783
+  C1=0.00000000000471
+  C2=0.00000000000684
+  RS1=504
+  RS2=500
+  RS3=545
+  RS4=11862
+  RS5=676
+  R2=11
.ends L_744824433_3.3m
****
.subckt L_744824220_20m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000077
+  DL4=0.000000485
+  DC3=0.000000000028
+  DC4=0.000000000011
+  DR3=17
+  dR4=50k
+  DR5=30
+  dR6=5k
+  Rdc=175.322m
+  ck=5pF
+  L1=18.2m
+  L2=0.7m
+  L3=23u
+  L4=4u
+  L5=2.2u
+  C1=32p
+  C2=23p
+  Rs1=46k
+  Rs2=39k
+  RS3=500
+  RS4=600
+  RS5=3000
+  R2=10.41
.ends L_744824220_20m
****
.subckt L_744824310_10m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=0.00975054658861754
+  L2=1.14140874719913E-06
+  L3=0.0000194215546747162
+  L4=1.85397202790917E-06
+  L5=1.37528846983612E-06
+  C1=1.06648809782419E-11
+  C2=1.54875317445924E-11
+  RS1=68798.4459196234
+  RS2=49005.5273080916
+  RS3=4486.62345566418
+  RS4=361.356712407375
+  RS5=1960.56329938029
+  R2=11.2784542155485
+  DL3=3.33880176803062E-06
+  DC3=1.51444689487349E-11
+  DL4=4.03878815013849E-09
+  DC4=6.73761021204444E-12
+  DR3=0.717429786820428
+  DR4=17180.6679766708
+  DR5=55.0109730646157
+  DR6=3197.74941444441
+  Rdc=85.225m
+  ck=4pF
.ends L_744824310_10m
****
.subckt XL_7448251201_1m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000003
+  DC3=0.00000000001
+  DL4=0.00000000951
+  DC4=0.00000000000463
+  DR3=0.18
+  DR4=2680
+  DR5=0.78
+  DR6=366
+  Rdc=5.598m
+  ck=5pF
+  L1=0.00022
+  L2=0.00019
+  L3=0.00022
+  L4=0.00064
+  L5=0.00000001398
+  C1=0.00000000000335
+  C2=0.00000000000531
+  RS1=560
+  RS2=550
+  RS3=1500
+  RS4=798
+  RS5=269
+  R2=7
.ends XL_7448251201_1m
****
.subckt XL_7448258022_2.2m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.00000058
+  DL4=0.000000025
+  DC3=0.0000000000165
+  DC4=0.00000000001
+  DR3=17
+  dR4=7k
+  DR5=23
+  dR6=3k
+  Rdc=11.1m
+  ck=1pF
+  L1=1.8m
+  L2=80u
+  L3=23u
+  L4=4u
+  L5=135n
+  C1=4.5p
+  C2=1.5p
+  RS1=4000
+  RS2=1600
+  RS3=1500
+  RS4=200
+  RS5=800
+  R2=1
.ends XL_7448258022_2.2m
****
.subckt XL_7448256033_3.3m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.00000085
+  DL4=0.000000058
+  DC3=0.0000000000144
+  DC4=0.000000000001
+  DR3=17
+  dR4=9k
+  DR5=23
+  dR6=2k
+  Rdc=18.752m
+  ck=4pF
+  L1=2.6m
+  L2=700u
+  L3=23u
+  L4=4u
+  L5=110.4n
+  C1=5p
+  C2=2.8p
+  Rs1=16k
+  Rs2=6k
+  RS3=500
+  RS4=600
+  RS5=900
+  R2=10.41
.ends XL_7448256033_3.3m
****
.subckt XL_744825605_5m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.00000133
+  DC3=0.00000000001775
+  DL4=0.00000003977
+  DC4=0.00000000002487
+  DR3=13
+  DR4=7090
+  DR5=13
+  DR6=6762
+  Rdc=35.042m
+  ck=2pF
+  L1=0.00034616
+  L2=0.00025028
+  L3=0.00025626
+  L4=0.00065136
+  L5=0.0000001087
+  C1=0.00000000000515
+  C2=0.00000000000874
+  RS1=2558
+  RS2=2548
+  RS3=6527
+  RS4=2609
+  RS5=674
+  R2=15
.ends XL_744825605_5m
****
.subckt XL_744825510_10m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000027
+  DL4=0.000000081
+  DC3=0.000000000037
+  DC4=0.000000000005
+  DR3=17
+  dR4=30k
+  DR5=23
+  dR6=12k
+  Rdc=40.604m
+  ck=5pF
+  L1=8m
+  L2=1m
+  L3=23u
+  L4=4u
+  L5=600.4n
+  C1=22p
+  C2=16p
+  Rs1=60k
+  RS2=6000
+  RS3=500
+  RS4=600
+  RS5=1600
+  R2=1.41
.ends XL_744825510_10m
****
.subckt XL_744825320_20m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.0000059
+  DL4=0.00000014
+  DC3=0.000000000036
+  DC4=0.000000000046
+  DR3=17
+  dR4=35k
+  DR5=23
+  dR6=9k
+  Rdc=123.197m
+  ck=5pF
+  L1=16m
+  L2=580u
+  L3=23u
+  L4=4u
+  L5=900.4n
+  C1=31p
+  C2=48p
+  Rs1=62k
+  Rs2=6k
+  RS3=500
+  RS4=600
+  RS5=1600
+  R2=1.41
.ends XL_744825320_20m
****
.subckt XL_744825433_33m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=0.0282615082580083
+  L2=0.00151069974592023
+  L3=0.0000635319123130355
+  L4=0.0000802861920160678
+  L5=8.4783967316618E-07
+  C1=3.31973088954225E-11
+  C2=8.99664633755108E-11
+  RS1=271189.203553144
+  RS2=68603.4021105262
+  RS3=958.938477130436
+  RS4=557.325344506158
+  RS5=1527.4005919289
+  R2=54.5016446977904
+  DL3=9.83880176803062E-06
+  DC3=4.9444689487349E-11
+  DL4=2.00387881501384E-07
+  DC4=4.17376102120444E-11
+  DR3=0.217429786820428
+  DR4=19180.6679766708
+  DR5=39.0109730646157
+  DR6=5197.74941444441
+  Rdc=187.34m
+  ck=4pF
.ends XL_744825433_33m
****
.subckt XXL_7448262510_1m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=0.00030889
+  L2=0.00039029
+  L3=0.00005
+  L4=0.00005
+  L5=0.00032526
+  C1=0.0000000000218
+  C2=0.00000000000527
+  RS1=3140
+  RS2=2206
+  RS3=3254
+  RS4=4188
+  RS5=3190
+  R2=0.054
+  DL3=0.00000049
+  DC3=0.0000000000129
+  DL4=0.00000003711
+  DC4=0.00000000000007
+  DR3=0.48
+  DR4=3680
+  DR5=18
+  DR6=366
+  Rdc=3.427m
+  ck=4pF
.ends XXL_7448262510_1m
****
.subckt XXL_7448261418_1.8m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=0.00140889
+  L2=0.00039029
+  L3=0.00005
+  L4=0.00005
+  L5=0.00012526
+  C1=0.0000000000098
+  C2=0.00000000000987
+  RS1=8140
+  RS2=8206
+  RS3=3254
+  RS4=4188
+  RS5=2500
+  R2=0.054
+  DL3=0.00000094
+  DC3=0.0000000000176
+  DL4=0.00000005111
+  DC4=0.00000000000233
+  DR3=0.48
+  DR4=6680
+  DR5=0.58
+  DR6=566
+  Rdc=7.79m
+  ck=4pF
.ends XXL_7448261418_1.8m
****
.subckt XXL_7448262013_1.3m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=0.00060889
+  L2=0.00059029
+  L3=0.00005
+  L4=0.00001
+  L5=0.00012526
+  C1=0.0000000000108
+  C2=0.00000000000687
+  RS1=4140
+  RS2=2206
+  RS3=2254
+  RS4=3188
+  RS5=2100
+  R2=0.054
+  DL3=0.00000062
+  DC3=0.0000000000148
+  DL4=0.00000003811
+  DC4=0.00000000000213
+  DR3=0.48
+  DR4=4680
+  DR5=0.58
+  DR6=446
+  Rdc=4.8m
+  ck=4pF
.ends XXL_7448262013_1.3m
****
.subckt XXL_7448263505_0.5m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  L1=0.000209496782810346
+  L2=0.000207729580657503
+  L3=0.000244939980673891
+  L4=4.35416881861321E-06
+  L5=0.0000181955270659663
+  C1=7.22232517664312E-11
+  C2=6.74966861088266E-11
+  RS1=12.914504794244
+  RS2=2355.13991346187
+  RS3=1395.50992687538
+  RS4=13415.8487785026
+  RS5=260.107405675112
+  R2=40.2708746893173
+  DL3=0.00000023
+  DC3=0.0000000000106
+  DL4=0.00000001211
+  DC4=0.00000000000033
+  DR3=0.48
+  DR4=1580
+  DR5=0.58
+  DR6=166
+  Rdc=1.84m
+  ck=4pF
.ends XXL_7448263505_0.5m
****
.subckt S_744822222_2.2m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.68u
+  DL4=3n
+  DC3=8.3p
+  DC4=2p
+  DR3=17
+  dR4=6k
+  DR5=30
+  dR6=2k
+  Rdc=0.079
+  ck=3pF
+  L1=1.75m
+  L2=0.58m
+  L3=23u
+  L4=4u
+  L5=210.4n
+  C1=6.5p
+  C2=8p
+  Rs1=17.5k
+  Rs2=6k
+  RS3=500
+  RS4=200
+  RS5=1200
+  R2=1.41
.ends S_744822222_2.2m
****
.subckt L_744824407_7m 1 2 3 4
X1  1  2  3  4  CMB  PARAMS:
+  DL3=0.00000228242
+  DC3=0.00000000001367
+  DL4=0.000000159
+  DC4=0.00000000000971
+  DR3=0.02
+  DR4=8278
+  DR5=28
+  DR6=821
+  Rdc=16.345m
+  ck=2pF
+  L1=0.00000897
+  L2=0.00016374
+  L3=0.00221744
+  L4=0.00443191
+  L5=0.00000010639
+  C1=0.00000000002399
+  C2=0.00000000001211
+  RS1=10
+  RS2=943
+  RS3=30928
+  RS4=30391
+  RS5=765
+  R2=4
.ends L_744824407_7m
****
.subckt L_744824801_1m  1 2 3 4
X1  1  2  3  4  CMB1  PARAMS:
+ L3=1150u
+ Rs3=6.4k
+ C1=12p
+ R2=1
+ L1=0.1p
+ Rs2=700
+ C2=0.1u
+ Rs1=10
+ L2=1u
+ L4=0.01u
+ Rs4=1
+ L5=0.01p
+ Rs5=0.1k
+ dR5=1
+ Rdc=1m
+ ck=3p
+ dR3=1k
+ dR6=2.8k
+ dR4=1k
+ dC3=2.1p
+ dL3=0.2u
+ dC4=1p
+ dL4=0.245u
.ends
****
.subckt XL_744825410_10m  1 2 3 4
X1  1  2  3  4  CMB1  PARAMS:
+ L3=10m
+ Rs3=116.4k
+ C1=32p
+ R2=1
+ L1=0.1p
+ Rs2=700
+ C2=0.1u
+ Rs1=10
+ L2=1u
+ L4=0.01u
+ Rs4=1
+ L5=0.01p
+ Rs5=0.1k
+ dR5=1
+ Rdc=1m
+ ck=8p
+ dR3=1.1k
+ dR6=10.1k
+ dR4=1.1k
+ dC3=10.1p
+ dL3=0.30u
+ dC4=1p
+ dL4=2.4u
.ends
****
.subckt L_744824405_5m  1 2 3 4
X1  1  2  3  4  CMB1  PARAMS:
+ L3=5.6m
+ Rs3=44.0k
+ C1=14.5p
+ R2=1
+ L1=0.1p
+ Rs2=100
+ C2=0.1u
+ Rs1=10
+ L2=1u
+ L4=0.01u
+ Rs4=1
+ L5=0.01p
+ Rs5=0.01k
+ dR5=1
+ Rdc=1m
+ ck=5p
+ dR3=2.1k
+ dR6=23.4k
+ dR4=1.1k
+ dC3=10p
+ dL3=0.60u
+ dC4=0.8p
+ dL4=1.0u
.ends