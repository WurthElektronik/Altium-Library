**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT High Current Flat Wire Inductor 
* Matchcode:             WE-HCM
* Library Type:          spice
* Version:               rev
* Created/modified by:   Ella
* Date and Time:         7/25/2023
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
.subckt 1050_744303012_0.12u 1 2
Rp 1 2 71.54
Cp 1 2 11p
Rs 1 N3 0.000325
L1 N3 2 0.12144u
.ends 1050_744303012_0.12u
*******
.subckt 1050_744303015_0.155u 1 2
Rp 1 2 69.77
Cp 1 2 20.21p
Rs 1 N3 0.000325
L1 N3 2 0.1706u
.ends 1050_744303015_0.155u
*******
.subckt 1050_744303022_0.22u 1 2
Rp 1 2 84.88
Cp 1 2 18.52p
Rs 1 N3 0.000325
L1 N3 2 0.26084u
.ends 1050_744303022_0.22u
*******
.subckt 1052_744306020_0.2u 1 2
Rp 1 2 53.9
Cp 1 2 34.0207585052126p
Rs 1 N3 0.00026
L1 N3 2 0.22133u
.ends 1052_744306020_0.2u
*******
.subckt 1052_744306025_0.25u 1 2
Rp 1 2 55.47
Cp 1 2 53.8437526344042p
Rs 1 N3 0.00026
L1 N3 2 0.32579u
.ends 1052_744306025_0.25u
*******
.subckt 1052_744306030_0.3u 1 2
Rp 1 2 53.22
Cp 1 2 71.8365539553462p
Rs 1 N3 0.00026
L1 N3 2 0.36692u
.ends 1052_744306030_0.3u
*******
.subckt 1070_744308015_0.15u 1 2
Rp 1 2 57.41
Cp 1 2 35.5686649908743p
Rs 1 N3 0.00037
L1 N3 2 0.19782u
.ends 1070_744308015_0.15u
*******
.subckt 1070_744308020_0.2u 1 2
Rp 1 2 61.66
Cp 1 2 58.2264493040575p
Rs 1 N3 0.00037
L1 N3 2 0.21483u
.ends 1070_744308020_0.2u
*******
.subckt 1070_744308025_0.25u 1 2
Rp 1 2 64.55
Cp 1 2 54.1116141235027p
Rs 1 N3 0.00037
L1 N3 2 0.29257u
.ends 1070_744308025_0.25u
*******
.subckt 1070_744308033_0.33u 1 2
Rp 1 2 69.73
Cp 1 2 53.0553512086678p
Rs 1 N3 0.00037
L1 N3 2 0.38974u
.ends 1070_744308033_0.33u
*******
.subckt 1070_744308040_0.4u 1 2
Rp 1 2 50.667
Cp 1 2 80.7876010519523p
Rs 1 N3 0.00037
L1 N3 2 0.501667u
.ends 1070_744308040_0.4u
*******
.subckt 1088_7443082010B_0.1u 1 2
Rp 1 2 29
Cp 1 2 46p
Rs 1 N3 0.000114
L1 N3 2 0.109u
.ends 1088_7443082010B_0.1u
*******
.subckt 1088_7443082012B_0.12u 1 2
Rp 1 2 31
Cp 1 2 56p
Rs 1 N3 0.000114
L1 N3 2 0.129u
.ends 1088_7443082012B_0.12u
*******
.subckt 1088_7443082015B_0.15u 1 2
Rp 1 2 32
Cp 1 2 63p
Rs 1 N3 0.000114
L1 N3 2 0.162u
.ends 1088_7443082015B_0.15u
*******
.subckt 1190_744301025_0.25u 1 2
Rp 1 2 45.7
Cp 1 2 1.44229442907223p
Rs 1 N3 0.00032
L1 N3 2 0.281u
.ends 1190_744301025_0.25u
*******
.subckt 1190_744301033_0.33u 1 2
Rp 1 2 34.58
Cp 1 2 6.74413480406324p
Rs 1 N3 0.00032
L1 N3 2 0.284u
.ends 1190_744301033_0.33u
*******
.subckt 1190_744301047_0.47u 1 2
Rp 1 2 47.76
Cp 1 2 4.30743392010698p
Rs 1 N3 0.00032
L1 N3 2 0.486u
.ends 1190_744301047_0.47u
*******
.subckt 1240_744304010_0.1u 1 2
Rp 1 2 41.01
Cp 1 2 21.5730752009037p
Rs 1 N3 0.00017
L1 N3 2 0.1065u
.ends 1240_744304010_0.1u
*******
.subckt 1240_744304016_0.16u 1 2
Rp 1 2 59.08
Cp 1 2 22.9840809293165p
Rs 1 N3 0.00017
L1 N3 2 0.1722u
.ends 1240_744304016_0.16u
*******
.subckt 1240_744304022_0.22u 1 2
Rp 1 2 51.23
Cp 1 2 23.1813818162177p
Rs 1 N3 0.00017
L1 N3 2 0.223u
.ends 1240_744304022_0.22u
*******
.subckt 1350_744305022_0.22u 1 2
Rp 1 2 55.28
Cp 1 2 88.8408246022065p
Rs 1 N3 0.000155
L1 N3 2 0.22u
.ends 1350_744305022_0.22u
*******
.subckt 1350_744305033_0.33u 1 2
Rp 1 2 58.24
Cp 1 2 143.928612643143p
Rs 1 N3 0.000155
L1 N3 2 0.36362u
.ends 1350_744305033_0.33u
*******
.subckt 1350_744305040_0.4u 1 2
Rp 1 2 62.85
Cp 1 2 131.044077014429p
Rs 1 N3 0.000155
L1 N3 2 0.48324u
.ends 1350_744305040_0.4u
*******
.subckt 1390_744309012_0.12u 1 2
Rp 1 2 32
Cp 1 2 56p
Rs 1 N3 0.000165
L1 N3 2 0.12u
.ends 1390_744309012_0.12u
*******
.subckt 1390_744309025_0.25u 1 2
Rp 1 2 35
Cp 1 2 76p
Rs 1 N3 0.000165
L1 N3 2 0.239u
.ends 1390_744309025_0.25u
*******
.subckt 1390_744309033_0.33u 1 2
Rp 1 2 38
Cp 1 2 96.43p
Rs 1 N3 0.000165
L1 N3 2 0.339u
.ends 1390_744309033_0.33u
*******
.subckt 1390_744309047_0.47u 1 2
Rp 1 2 39
Cp 1 2 120p
Rs 1 N3 0.000165
L1 N3 2 0.434u
.ends 1390_744309047_0.47u
*******
.subckt 1820_74431821100_1u 1 2
Rp 1 2 163.9
Cp 1 2 33.57p
Rs 1 N3 0.00033
L1 N3 2 0.7717u
.ends 1820_74431821100_1u
*******
.subckt 7050_744302007_0.072u 1 2
Rp 1 2 42.42
Cp 1 2 18.39p
Rs 1 N3 0.000235
L1 N3 2 0.077366u
.ends 7050_744302007_0.072u
*******
.subckt 7050_744302010_0.105u 1 2
Rp 1 2 35.46
Cp 1 2 50.45p
Rs 1 N3 0.000235
L1 N3 2 0.1178u
.ends 7050_744302010_0.105u
*******
.subckt 7050_744302015_0.15u 1 2
Rp 1 2 51.16
Cp 1 2 46.07p
Rs 1 N3 0.000235
L1 N3 2 0.16722u
.ends 7050_744302015_0.15u
*******
.subckt 7070_744307012_0.12u 1 2
Rp 1 2 41.79
Cp 1 2 35.4705123346616p
Rs 1 N3 0.00029
L1 N3 2 0.16394u
.ends 7070_744307012_0.12u
*******
.subckt 7070_744307016_0.16u 1 2
Rp 1 2 42.31
Cp 1 2 53.4563594187636p
Rs 1 N3 0.00029
L1 N3 2 0.18954u
.ends 7070_744307016_0.16u
*******
.subckt 7070_744307022_0.22u 1 2
Rp 1 2 36
Cp 1 2 78.376p
Rs 1 N3 0.00029
L1 N3 2 0.228u
.ends 7070_744307022_0.22u
*******
.subckt 1012_74431012007_0.07u 1 2
Rp 1 2 38.094
Cp 1 2 15.977p
Rs 1 N3 0.000125
L1 N3 2 0.071251u
.ends 1012_74431012007_0.07u
*******
.subckt 1012_74431012010_0.1u 1 2
Rp 1 2 33.974
Cp 1 2 35.541p
Rs 1 N3 0.000125
L1 N3 2 0.099838u
.ends 1012_74431012010_0.1u
*******
.subckt 1012_74431012012_0.12u 1 2
Rp 1 2 35.911
Cp 1 2 36.528p
Rs 1 N3 0.000125
L1 N3 2 0.12274u
.ends 1012_74431012012_0.12u
*******
.subckt 1012_74431012015_0.15u 1 2
Rp 1 2 41.646
Cp 1 2 33.261p
Rs 1 N3 0.000125
L1 N3 2 0.151517u
.ends 1012_74431012015_0.15u
*******
.subckt 1078_7443081010_0.1u 1 2
Rp 1 2 36.968
Cp 1 2 39.578587360283p
Rs 1 N3 0.00029
L1 N3 2 0.1u
.ends 1078_7443081010_0.1u
*******
.subckt 1078_7443081012_0.12u 1 2
Rp 1 2 36.968
Cp 1 2 38.5474432532583p
Rs 1 N3 0.00029
L1 N3 2 0.12u
.ends 1078_7443081012_0.12u
*******
.subckt 1078_7443081015_0.15u 1 2
Rp 1 2 37.033
Cp 1 2 38.3077284683456p
Rs 1 N3 0.00029
L1 N3 2 0.143u
.ends 1078_7443081015_0.15u
*******
.subckt 1078_7443081018_0.18u 1 2
Rp 1 2 38.971
Cp 1 2 52.042849914902p
Rs 1 N3 0.00029
L1 N3 2 0.18u
.ends 1078_7443081018_0.18u
*******
.subckt 1078_7443081022_0.22u 1 2
Rp 1 2 42.567
Cp 1 2 62.2702588882962p
Rs 1 N3 0.00029
L1 N3 2 0.22u
.ends 1078_7443081022_0.22u
*******
.subckt 1078_7443081030_0.3u 1 2
Rp 1 2 43.708
Cp 1 2 77.5338105619256p
Rs 1 N3 0.00029
L1 N3 2 0.3u
.ends 1078_7443081030_0.3u
*******
.subckt 1078_7443081040_0.4u 1 2
Rp 1 2 48.258
Cp 1 2 86.8665840554908p
Rs 1 N3 0.00029
L1 N3 2 0.4u
.ends 1078_7443081040_0.4u
*******
.subckt 1088_7443082010_0.1u 1 2
Rp 1 2 30.8
Cp 1 2 28.6099325913374p
Rs 1 N3 0.00018
L1 N3 2 0.1002u
.ends 1088_7443082010_0.1u
*******
.subckt 1088_7443082012_0.12u 1 2
Rp 1 2 38.47
Cp 1 2 43.1686692694493p
Rs 1 N3 0.00018
L1 N3 2 0.11975u
.ends 1088_7443082012_0.12u
*******
.subckt 1088_7443082015A_0.15u 1 2
Rp 1 2 33.62
Cp 1 2 54.9212125286487p
Rs 1 N3 0.00015
L1 N3 2 0.14707u
.ends 1088_7443082015A_0.15u
*******
.subckt 1088_7443082015_0.15u 1 2
Rp 1 2 31.74
Cp 1 2 45.6283316431974p
Rs 1 N3 0.00018
L1 N3 2 0.13987u
.ends 1088_7443082015_0.15u
*******
.subckt 1088_7443082017_0.17u 1 2
Rp 1 2 30
Cp 1 2 45.7790904930195p
Rs 1 N3 0.00018
L1 N3 2 0.17644u
.ends 1088_7443082017_0.17u
*******
.subckt 1088_7443082018A_0.18u 1 2
Rp 1 2 36.81
Cp 1 2 63.2375281674737p
Rs 1 N3 0.00015
L1 N3 2 0.18133u
.ends 1088_7443082018A_0.18u
*******
.subckt 1088_7443082018_0.18u 1 2
Rp 1 2 30.33
Cp 1 2 50.2370433090238p
Rs 1 N3 0.00018
L1 N3 2 0.1795u
.ends 1088_7443082018_0.18u
*******
.subckt 1088_7443082022_0.22u 1 2
Rp 1 2 33.66
Cp 1 2 43.5991482113114p
Rs 1 N3 0.00018
L1 N3 2 0.21486u
.ends 1088_7443082022_0.22u
*******
.subckt 1323_74431323012_0.12u 1 2
Rp 1 2 67.84
Cp 1 2 14.6905656182035p
Rs 1 N3 0.0007
L1 N3 2 0.11974u
.ends 1323_74431323012_0.12u
*******
.subckt 1323_74431323016_0.16u 1 2
Rp 1 2 66.58
Cp 1 2 12.2999362792959p
Rs 1 N3 0.0007
L1 N3 2 0.16128u
.ends 1323_74431323016_0.16u
*******
.subckt 1411_7443091062_0.62u 1 2
Rp 1 2 59
Cp 1 2 69p
Rs 1 N3 0.00042
L1 N3 2 0.598u
.ends 1411_7443091062_0.62u
*******
.subckt 1411_7443091080_0.8u 1 2
Rp 1 2 79
Cp 1 2 96p
Rs 1 N3 0.00042
L1 N3 2 0.767u
.ends 1411_7443091080_0.8u
*******
.subckt 1411_7443091100_1u 1 2
Rp 1 2 103
Cp 1 2 57p
Rs 1 N3 0.00042
L1 N3 2 1u
.ends 1411_7443091100_1u
*******
.subckt 1411_7443091120_1.2u 1 2
Rp 1 2 104
Cp 1 2 104p
Rs 1 N3 0.00042
L1 N3 2 1.2u
.ends 1411_7443091120_1.2u
*******
.subckt 1411_7443091150_1.5u 1 2
Rp 1 2 107
Cp 1 2 93p
Rs 1 N3 0.00042
L1 N3 2 1.5u
.ends 1411_7443091150_1.5u
*******
.subckt 1435_74431435010_0.1u 1 2
Rp 1 2 48
Cp 1 2 31.5715491822168p
Rs 1 N3 0.00028
L1 N3 2 0.106u
.ends 1435_74431435010_0.1u
*******
.subckt 1435_74431435012_0.12u 1 2
Rp 1 2 51
Cp 1 2 26.1636067867387p
Rs 1 N3 0.00028
L1 N3 2 0.134u
.ends 1435_74431435012_0.12u
*******
.subckt 1435_74431435015_0.15u 1 2
Rp 1 2 46
Cp 1 2 24.2560442239891p
Rs 1 N3 0.00028
L1 N3 2 0.148u
.ends 1435_74431435015_0.15u
*******
.subckt 1435_74431435018_0.18u 1 2
Rp 1 2 52
Cp 1 2 32.232498721889p
Rs 1 N3 0.00028
L1 N3 2 0.198u
.ends 1435_74431435018_0.18u
*******
.subckt 1435_74431435022_0.22u 1 2
Rp 1 2 52
Cp 1 2 31.4115772700659p
Rs 1 N3 0.00028
L1 N3 2 0.224u
.ends 1435_74431435022_0.22u
*******
.subckt 4030_744340300025_0.025u 1 2
Rp 1 2 38.094
Cp 1 2 15.977p
Rs 1 N3 0.00027
L1 N3 2 0.071251u
.ends 4030_744340300025_0.025u
*******
.subckt 4030_744340300030_0.03u 1 2
Rp 1 2 33.974
Cp 1 2 35.541p
Rs 1 N3 0.00027
L1 N3 2 0.099838u
.ends 4030_744340300030_0.03u
*******
.subckt 4030_744340300055_0.055u 1 2
Rp 1 2 35.911
Cp 1 2 36.528p
Rs 1 N3 0.00027
L1 N3 2 0.12274u
.ends 4030_744340300055_0.055u
*******
.subckt 4030_744340300075_0.075u 1 2
Rp 1 2 41.646
Cp 1 2 33.261p
Rs 1 N3 0.00027
L1 N3 2 0.151517u
.ends 4030_744340300075_0.075u
*******
.subckt 4035_74434035007_0.07u 1 2
Rp 1 2 26.693
Cp 1 2 51.328p
Rs 1 N3 0.00038
L1 N3 2 0.069034u
.ends 4035_74434035007_0.07u
*******
.subckt 4035_74434035010_0.1u 1 2
Rp 1 2 31.361
Cp 1 2 58.945p
Rs 1 N3 0.00038
L1 N3 2 0.08884u
.ends 4035_74434035010_0.1u
*******
.subckt 5030_74435030010_0.1u 1 2
Rp 1 2 37.557
Cp 1 2 37.678p
Rs 1 N3 0.00031
L1 N3 2 0.096909u
.ends 5030_74435030010_0.1u
*******
.subckt 9065_744300006_0.06u 1 2
Rp 1 2 27.774
Cp 1 2 26.65p
Rs 1 N3 0.00022
L1 N3 2 0.061889u
.ends 9065_744300006_0.06u
*******
.subckt 9065_744300008_0.08u 1 2
Rp 1 2 28.724
Cp 1 2 36.05p
Rs 1 N3 0.00022
L1 N3 2 0.078758u
.ends 9065_744300008_0.08u
*******
.subckt 9065_744300010_0.1u 1 2
Rp 1 2 30.193
Cp 1 2 46.623p
Rs 1 N3 0.00022
L1 N3 2 0.098291u
.ends 9065_744300010_0.1u
*******
.subckt 9065_744300015_0.15u 1 2
Rp 1 2 33.62
Cp 1 2 67.437p
Rs 1 N3 0.00022
L1 N3 2 0.146178u
.ends 9065_744300015_0.15u
*******
.subckt 9065_744300022_0.22u 1 2
Rp 1 2 34.612
Cp 1 2 80.172p
Rs 1 N3 0.00022
L1 N3 2 0.218406u
.ends 9065_744300022_0.22u
*******
