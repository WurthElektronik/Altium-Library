**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Universal Offline Standard Transformers
* Matchcode:              WE-UOST
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Toby      
* Date and Time:          2022-05-17
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************

.subckt 760875532		9  7  12  11  1  2  3  5		
.param RxLkg=14868.88ohm					
.param Leakage=49uh					
Rlkg	9	9a	{RxLkg}		
L_Lkg	9	9a	{Leakage}	Rser=0.01mohm	
Lpri1	9a	7	1451uH	Rser=5500mohm	
Laux1	12	11	15uH	Rser=300mohm	
Lsec1	1	2	5.859uH	Rser=70mohm	
Lsec2	3	5	2.871uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=18.1pf					
.param Rdmp1=455169.65ohm					
Cpri1	9	7	{Cprm1}	Rser=10mohm	
Rdmp1	9	7	{Rdmp1}		
Rg3	9	0	20meg		
Rg5	12	0	20meg		
Rg7	7	0	20meg		
Rg9	11	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	2	0	20meg		
Rg20	5	0	20meg		
.ends					

.subckt 760875131		9  7  12  11  1  4  3  6		
.param RxLkg=15989.98ohm					
.param Leakage=45uh					
Rlkg	9	9a	{RxLkg}		
L_Lkg	9	9a	{Leakage}	Rser=0.01mohm	
Lpri1	9a	7	1455uH	Rser=3400mohm	
Laux1	12	11	15uH	Rser=280mohm	
Lsec1	1	4	11.484uH	Rser=110mohm	
Lsec2	3	6	11.484uH	Rser=110mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=13.2pf					
.param Rdmp1=532999.47ohm					
Cpri1	9	7	{Cprm1}	Rser=10mohm	
Rdmp1	9	7	{Rdmp1}		
Rg3	9	0	20meg		
Rg5	12	0	20meg		
Rg7	7	0	20meg		
Rg9	11	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	4	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt 760875112		9  7  12  11  1  4  3  6		
.param RxLkg=13820.44ohm					
.param Leakage=38uh					
Rlkg	9	9a	{RxLkg}		
L_Lkg	9	9a	{Leakage}	Rser=0.01mohm	
Lpri1	9a	7	1462uH	Rser=3400mohm	
Laux1	12	11	18.984uH	Rser=300mohm	
Lsec1	1	4	2.871uH	Rser=20mohm	
Lsec2	3	6	2.871uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=12.6pf					
.param Rdmp1=545543.85ohm					
Cpri1	9	7	{Cprm1}	Rser=10mohm	
Rdmp1	9	7	{Rdmp1}		
Rg3	9	0	20meg		
Rg5	12	0	20meg		
Rg7	7	0	20meg		
Rg9	11	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	4	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt 760871142		9  7  12  11  1  4  3  6		
.param RxLkg=13403.39ohm					
.param Leakage=32uh					
Rlkg	9	9a	{RxLkg}		
L_Lkg	9	9a	{Leakage}	Rser=0.01mohm	
Lpri1	9a	7	1218uH	Rser=2400mohm	
Laux1	12	11	16.327uH	Rser=300mohm	
Lsec1	1	4	46.492uH	Rser=430mohm	
Lsec2	3	6	46.492uH	Rser=460mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=11.4pf					
.param Rdmp1=523569.98ohm					
Cpri1	9	7	{Cprm1}	Rser=10mohm	
Rdmp1	9	7	{Rdmp1}		
Rg3	9	0	20meg		
Rg5	12	0	20meg		
Rg7	7	0	20meg		
Rg9	11	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	4	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt 760871534		9  7  12  11  1  2  3  5		
.param RxLkg=10527.1ohm					
.param Leakage=26uh					
Rlkg	9	9a	{RxLkg}		
L_Lkg	9	9a	{Leakage}	Rser=0.01mohm	
Lpri1	9a	7	1224uH	Rser=2400mohm	
Laux1	12	11	20.663uH	Rser=300mohm	
Lsec1	1	2	5.166uH	Rser=200mohm	
Lsec2	3	5	3.125uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=12.2pf					
.param Rdmp1=506110.58ohm					
Cpri1	9	7	{Cprm1}	Rser=10mohm	
Rdmp1	9	7	{Rdmp1}		
Rg3	9	0	20meg		
Rg5	12	0	20meg		
Rg7	7	0	20meg		
Rg9	11	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	2	0	20meg		
Rg20	5	0	20meg		
.ends					

.subckt 760871543		9  7  12  11  1  2  3  5		
.param RxLkg=12729.29ohm					
.param Leakage=30uh					
Rlkg	9	9a	{RxLkg}		
L_Lkg	9	9a	{Leakage}	Rser=0.01mohm	
Lpri1	9a	7	1280uH	Rser=2400mohm	
Laux1	12	11	17.11uH	Rser=200mohm	
Lsec1	1	2	32.349uH	Rser=400mohm	
Lsec2	3	5	2.406uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=10.6pf					
.param Rdmp1=555845.82ohm					
Cpri1	9	7	{Cprm1}	Rser=10mohm	
Rdmp1	9	7	{Rdmp1}		
Rg3	9	0	20meg		
Rg5	12	0	20meg		
Rg7	7	0	20meg		
Rg9	11	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	2	0	20meg		
Rg20	5	0	20meg		
.ends					

.subckt 760871113		9  7  12  11  1  4  3  6		
.param RxLkg=12013.76ohm					
.param Leakage=30uh					
Rlkg	9	9a	{RxLkg}		
L_Lkg	9	9a	{Leakage}	Rser=0.01mohm	
Lpri1	9a	7	1280uH	Rser=2400mohm	
Laux1	12	11	17.11uH	Rser=300mohm	
Lsec1	1	4	2.406uH	Rser=20mohm	
Lsec2	3	6	2.406uH	Rser=20mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=11.9pf					
.param Rdmp1=524601.05ohm					
Cpri1	9	7	{Cprm1}	Rser=10mohm	
Rdmp1	9	7	{Rdmp1}		
Rg3	9	0	20meg		
Rg5	12	0	20meg		
Rg7	7	0	20meg		
Rg9	11	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	4	0	20meg		
Rg20	6	0	20meg		
.ends					

.subckt 760871135		9  7  12  11  1  4  3  6		
.param RxLkg=19686.23ohm					
.param Leakage=47uh					
Rlkg	9	9a	{RxLkg}		
L_Lkg	9	9a	{Leakage}	Rser=0.01mohm	
Lpri1	9a	7	1203uH	Rser=2400mohm	
Laux1	12	11	15.206uH	Rser=400mohm	
Lsec1	1	4	11.421uH	Rser=80mohm	
Lsec2	3	6	11.421uH	Rser=80mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=11.4pf					
.param Rdmp1=523569.98ohm					
Cpri1	9	7	{Cprm1}	Rser=10mohm	
Rdmp1	9	7	{Rdmp1}		
Rg3	9	0	20meg		
Rg5	12	0	20meg		
Rg7	7	0	20meg		
Rg9	11	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	4	0	20meg		
Rg20	6	0	20meg		
.ends					
