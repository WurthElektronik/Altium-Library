**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  Aluminum Electrolytic Capacitors
* Matchcode:              WCAP-AIG5
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          9/9/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 861021483001_33uF 1 2
Rser 1 3 0.322
Lser 2 4 1.3338018891E-08
C1 3 4 0.000033
Rpar 3 4 1515151.51515152
.ends 861021483001_33uF
*******
.subckt 861021483002_47uF 1 2
Rser 1 3 0.543
Lser 2 4 1.379797903E-08
C1 3 4 0.000047
Rpar 3 4 1063829.78723404
.ends 861021483002_47uF
*******
.subckt 861021483003_56uF 1 2
Rser 1 3 0.499
Lser 2 4 1.5328561293E-08
C1 3 4 0.000056
Rpar 3 4 892857.142857143
.ends 861021483003_56uF
*******
.subckt 861021483004_68uF 1 2
Rser 1 3 0.357
Lser 2 4 1.2697542772E-08
C1 3 4 0.000068
Rpar 3 4 735294.117647059
.ends 861021483004_68uF
*******
.subckt 861021483005_82uF 1 2
Rser 1 3 0.312
Lser 2 4 1.400840076E-08
C1 3 4 0.000082
Rpar 3 4 609756.097560976
.ends 861021483005_82uF
*******
.subckt 861021483006_100uF 1 2
Rser 1 3 0.264
Lser 2 4 1.3254828961E-08
C1 3 4 0.0001
Rpar 3 4 500000
.ends 861021483006_100uF
*******
.subckt 861021483007_120uF 1 2
Rser 1 3 0.221
Lser 2 4 1.3231589496E-08
C1 3 4 0.00012
Rpar 3 4 416666.666666667
.ends 861021483007_120uF
*******
.subckt 861021483008_150uF 1 2
Rser 1 3 0.182
Lser 2 4 1.2737604723E-08
C1 3 4 0.00015
Rpar 3 4 333333.333333333
.ends 861021483008_150uF
*******
.subckt 861021084013_470uF 1 2
Rser 1 3 0.15412
Lser 2 4 1.6735137504E-08
C1 3 4 0.00047
Rpar 3 4 106382.978723404
.ends 861021084013_470uF
*******
.subckt 861021484009_47uF 1 2
Rser 1 3 0.28
Lser 2 4 1.5516609918E-08
C1 3 4 0.000047
Rpar 3 4 1063829.78723404
.ends 861021484009_47uF
*******
.subckt 861021484010_56uF 1 2
Rser 1 3 0.432
Lser 2 4 1.4387829374E-08
C1 3 4 0.000056
Rpar 3 4 892857.142857143
.ends 861021484010_56uF
*******
.subckt 861021484011_68uF 1 2
Rser 1 3 0.353
Lser 2 4 1.5984962666E-08
C1 3 4 0.000068
Rpar 3 4 735294.117647059
.ends 861021484011_68uF
*******
.subckt 861021484012_82uF 1 2
Rser 1 3 0.323
Lser 2 4 1.6450787796E-08
C1 3 4 0.000082
Rpar 3 4 609756.097560976
.ends 861021484012_82uF
*******
.subckt 861021484013_100uF 1 2
Rser 1 3 0.285
Lser 2 4 1.80700838462865E-08
C1 3 4 0.0001
Rpar 3 4 500000
.ends 861021484013_100uF
*******
.subckt 861021484014_120uF 1 2
Rser 1 3 0.241
Lser 2 4 1.3748903207E-08
C1 3 4 0.00012
Rpar 3 4 416666.666666667
.ends 861021484014_120uF
*******
.subckt 861021484015_150uF 1 2
Rser 1 3 0.205
Lser 2 4 1.4130714112E-08
C1 3 4 0.00015
Rpar 3 4 333333.333333333
.ends 861021484015_150uF
*******
.subckt 861021484016_180uF 1 2
Rser 1 3 0.164
Lser 2 4 2.3322157863922E-08
C1 3 4 0.00018
Rpar 3 4 277777.777777778
.ends 861021484016_180uF
*******
.subckt 861021484017_220uF 1 2
Rser 1 3 0.153
Lser 2 4 1.4049168886E-08
C1 3 4 0.00022
Rpar 3 4 227272.727272727
.ends 861021484017_220uF
*******
.subckt 861021385017_220uF 1 2
Rser 1 3 0.27238
Lser 2 4 1.2413709855E-08
C1 3 4 0.00022
Rpar 3 4 227272.727272727
.ends 861021385017_220uF
*******
.subckt 861021485018_68uF 1 2
Rser 1 3 0.219
Lser 2 4 1.7567450756E-08
C1 3 4 0.000068
Rpar 3 4 735294.117647059
.ends 861021485018_68uF
*******
.subckt 861021485019_82uF 1 2
Rser 1 3 0.344
Lser 2 4 1.9515287897E-08
C1 3 4 0.000082
Rpar 3 4 609756.097560976
.ends 861021485019_82uF
*******
.subckt 861021085019_680uF 1 2
Rser 1 3 0.08259
Lser 2 4 1.9814528931E-08
C1 3 4 0.00068
Rpar 3 4 73529.4117647059
.ends 861021085019_680uF
*******
.subckt 861020785017_3.3mF 1 2
Rser 1 3 0.02898
Lser 2 4 1.879824471E-08
C1 3 4 0.0033
Rpar 3 4 15151.5151515152
.ends 861020785017_3.3mF
*******
.subckt 861021485020_100uF 1 2
Rser 1 3 0.265
Lser 2 4 1.6860174576E-08
C1 3 4 0.0001
Rpar 3 4 500000
.ends 861021485020_100uF
*******
.subckt 861021485021_120uF 1 2
Rser 1 3 0.224
Lser 2 4 1.549941039E-08
C1 3 4 0.00012
Rpar 3 4 416666.666666667
.ends 861021485021_120uF
*******
.subckt 861021485022_150uF 1 2
Rser 1 3 0.207
Lser 2 4 1.5123196725E-08
C1 3 4 0.00015
Rpar 3 4 333333.333333333
.ends 861021485022_150uF
*******
.subckt 861021485023_180uF 1 2
Rser 1 3 0.171
Lser 2 4 2.4651368900054E-08
C1 3 4 0.00018
Rpar 3 4 277777.777777778
.ends 861021485023_180uF
*******
.subckt 861021485024_220uF 1 2
Rser 1 3 0.156
Lser 2 4 1.5561763095E-08
C1 3 4 0.00022
Rpar 3 4 227272.727272727
.ends 861021485024_220uF
*******
.subckt 861021485025_270uF 1 2
Rser 1 3 0.116
Lser 2 4 1.03056721646618E-08
C1 3 4 0.00027
Rpar 3 4 185185.185185185
.ends 861021485025_270uF
*******
.subckt 861021485026_330uF 1 2
Rser 1 3 0.106
Lser 2 4 1.14239350877035E-08
C1 3 4 0.00033
Rpar 3 4 151515.151515152
.ends 861021485026_330uF
*******
.subckt 861021486027_150uF 1 2
Rser 1 3 0.219
Lser 2 4 1.7761290319E-08
C1 3 4 0.00015
Rpar 3 4 333333.333333333
.ends 861021486027_150uF
*******
.subckt 861021086027_1mF 1 2
Rser 1 3 0.089688
Lser 2 4 1.5452263797E-08
C1 3 4 0.001
Rpar 3 4 50000
.ends 861021086027_1mF
*******
.subckt 861020786024_4.7mF 1 2
Rser 1 3 0.024753
Lser 2 4 2.0343196996E-08
C1 3 4 0.0047
Rpar 3 4 10638.2978723404
.ends 861020786024_4.7mF
*******
.subckt 861021486028_180uF 1 2
Rser 1 3 0.182
Lser 2 4 1.16451389267057E-08
C1 3 4 0.00018
Rpar 3 4 277777.777777778
.ends 861021486028_180uF
*******
.subckt 861021386031_470uF 1 2
Rser 1 3 0.15642
Lser 2 4 1.3935747278E-08
C1 3 4 0.00047
Rpar 3 4 106382.978723404
.ends 861021386031_470uF
*******
.subckt 861021486029_220uF 1 2
Rser 1 3 0.153
Lser 2 4 2.7418263439451E-08
C1 3 4 0.00022
Rpar 3 4 227272.727272727
.ends 861021486029_220uF
*******
.subckt 861021486030_270uF 1 2
Rser 1 3 0.134
Lser 2 4 1.25222582623025E-08
C1 3 4 0.00027
Rpar 3 4 185185.185185185
.ends 861021486030_270uF
*******
.subckt 861020786030_10mF 1 2
Rser 1 3 0.028428
Lser 2 4 1.8963019704E-08
C1 3 4 0.01
Rpar 3 4 5000
.ends 861020786030_10mF
*******
.subckt 861021486031_330uF 1 2
Rser 1 3 0.125
Lser 2 4 2.69177695361617E-08
C1 3 4 0.00033
Rpar 3 4 151515.151515152
.ends 861021486031_330uF
*******
.subckt S861021486042_560uF 1 2
Rser 1 3 0.11
Lser 2 4 0.0000000096
C1 3 4 0.00056
Rpar 3 4 298804.780876494
.ends S861021486042_560uF
*******
.subckt 861021486032_390uF 1 2
Rser 1 3 0.109
Lser 2 4 2.80110841341855E-08
C1 3 4 0.00039
Rpar 3 4 128205.128205128
.ends 861021486032_390uF
*******
.subckt 861021386035_1mF 1 2
Rser 1 3 0.08386
Lser 2 4 1.4301110772E-08
C1 3 4 0.001
Rpar 3 4 50000
.ends 861021386035_1mF
*******
