**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT Wire Wound Ceramic Inductor
* Matchcode:             WE-KI
* Library Type:          LTspice
* Version:               rev21a
* Created/modified by:   Ella
* Date and Time:         5/24/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Wurth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Wurth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Wurth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Wurth Elektronik eiSos guarantee that the simulation model is current.
* Wurth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Wurth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0402_744765010A_1n 1 2
C1 1 N7 389.9518f
L1 1 N1 1n
L2 N1 N2 96.3426p
L3 N2 N3 139.4502p
L4 N3 N4 103.4194p
L5 N4 N5 63.1189p
L6 N5 N6 49.9792p
R1 2 N1 342.6049m
R2 2 N2 120.7838m
R3 2 N3 121.8758m
R4 2 N4 104.9031m
R5 2 N5 85.9424m
R6 2 N6 69.4743m
R7 2 N7 1.963
R8 2 1 1000000
.ends 0402_744765010A_1n
*******
.subckt 0402_744765019A_1.9n 1 2
C1 1 N7 268.5623f
L1 1 N1 1.7n
L2 N1 N2 205.5140p
L3 N2 N3 360.8888p
L4 N3 N4 330.0807p
L5 N4 N5 76.3595p
L6 N5 N6 54.0235p
R1 2 N1 365.6141m
R2 2 N2 363.8721m
R3 2 N3 329.5292m
R4 2 N4 271.9021m
R5 2 N5 245.0317m
R6 2 N6 90.3834m
R7 2 N7 1.9367
R8 2 1 1000000
.ends 0402_744765019A_1.9n
*******
.subckt 0402_744765020A_2n 1 2
C1 1 N7 0.3909p
L1 1 N1 1.8n
L2 N1 N2 113.5986p
L3 N2 N3 164.9783p
L4 N3 N4 127.9698p
L5 N4 N5 76.0574p
L6 N5 N6 53.8163p
R1 2 N1 408.3139m
R2 2 N2 156.8311m
R3 2 N3 143.0775m
R4 2 N4 122.8693m
R5 2 N5 103.3572m
R6 2 N6 89.5015m
R7 2 N7 1.9392
R8 2 1 1000000
.ends 0402_744765020A_2n
*******
.subckt 0402_744765022A_2.2n 1 2
C1 1 N7 0.35181p
L1 1 N1 2n
L2 N1 N2 134.6801p
L3 N2 N3 191.5544p
L4 N3 N4 209.2749p
L5 N4 N5 117.7200p
L6 N5 N6 65.4777p
R1 2 N1 423.9170m
R2 2 N2 244.3270m
R3 2 N3 218.5825m
R4 2 N4 184.8275m
R5 2 N5 161.4858m
R6 2 N6 152.4895m
R7 2 N7 1.9339
R8 2 1 1000000
.ends 0402_744765022A_2.2n
*******
.subckt 0402_744765024A_2.4n 1 2
C1 1 N7 295.2228f
L1 1 N1 2.2n
L2 N1 N2 134.4912p
L3 N2 N3 191.5524p
L4 N3 N4 209.5138p
L5 N4 N5 117.8466p
L6 N5 N6 65.5144p
R1 2 N1 538.3200m
R2 2 N2 217.2103m
R3 2 N3 218.7924m
R4 2 N4 185.0361m
R5 2 N5 161.6736m
R6 2 N6 152.6719m
R7 2 N7 1.9354
R8 2 1 1000000
.ends 0402_744765024A_2.4n
*******
.subckt 0402_744765027A_2.7n 1 2
C1 1 N7 212.4513f
L1 1 N1 2.5n
L2 N1 N2 145.0852p
L3 N2 N3 191.5524p
L4 N3 N4 212.7290p
L5 N4 N5 120.2424p
L6 N5 N6 66.1591p
R1 2 N1 724.8729m
R2 2 N2 356.5225m
R3 2 N3 222.8469m
R4 2 N4 188.9472m
R5 2 N5 165.1597m
R6 2 N6 156.0427m
R7 2 N7 1.931
R8 2 1 1000000
.ends 0402_744765027A_2.7n
*******
.subckt 0402_744765033A_3.3n 1 2
C1 1 N7 221.3170f
L1 1 N1 3.1n
L2 N1 N2 159.8447p
L3 N2 N3 191.5524p
L4 N3 N4 212.7290p
L5 N4 N5 132.5429p
L6 N5 N6 69.5011p
R1 2 N1 561.2163m
R2 2 N2 668.7847m
R3 2 N3 247.4353m
R4 2 N4 206.5131m
R5 2 N5 179.0585m
R6 2 N6 168.9615m
R7 2 N7 1.9286
R8 2 1 1000000
.ends 0402_744765033A_3.3n
*******
.subckt 0402_744765036A_3.6n 1 2
C1 1 N7 139.8032f
L1 1 N1 3.4n
L2 N1 N2 148.6566p
L3 N2 N3 191.8588p
L4 N3 N4 212.7290p
L5 N4 N5 137.7992p
L6 N5 N6 70.8751p
R1 2 N1 727.2652m
R2 2 N2 370.5498m
R3 2 N3 253.9939m
R4 2 N4 213.9650m
R5 2 N5 185.1919m
R6 2 N6 174.7227m
R7 2 N7 1.9207
R8 2 1 1000000
.ends 0402_744765036A_3.6n
*******
.subckt 0402_744765039A_3.9n 1 2
C1 1 N7 166.4000f
L1 1 N1 3.7n
L2 N1 N2 147.1866p
L3 N2 N3 191.8588p
L4 N3 N4 212.7290p
L5 N4 N5 139.6005p
L6 N5 N6 71.3408p
R1 2 N1 668.4030m
R2 2 N2 399.5452m
R3 2 N3 256.9274m
R4 2 N4 216.3665m
R5 2 N5 187.0541m
R6 2 N6 176.4355m
R7 2 N7 1.9211
R8 2 1 1000000
.ends 0402_744765039A_3.9n
*******
.subckt 0402_744765043A_4.3n 1 2
C1 1 N7 234.8940f
L1 1 N1 4n
L2 N1 N2 183.2147p
L3 N2 N3 191.8588p
L4 N3 N4 212.7290p
L5 N4 N5 254.3259p
L6 N5 N6 100.8976p
R1 2 N1 759.9111m
R2 2 N2 942.7394m
R3 2 N3 435.0905m
R4 2 N4 363.8248m
R5 2 N5 298.4430m
R6 2 N6 278.5925m
R7 2 N7 1.8927
R8 2 1 1000000
.ends 0402_744765043A_4.3n
*******
.subckt 0402_744765047A_4.7n 1 2
C1 1 N7 202.4121f
L1 1 N1 4.4n
L2 N1 N2 135.8640p
L3 N2 N3 131.1227p
L4 N3 N4 82.6537p
L5 N4 N5 47.1729p
L6 N5 N6 369.1065p
R1 2 N1 1.0836
R2 2 N2 1.2101
R3 2 N3 929.8133m
R4 2 N4 734.5717m
R5 2 N5 602.3623m
R6 2 N6 369.4921m
R7 2 N7 1.9766
R8 2 1 1000000
.ends 0402_744765047A_4.7n
*******
.subckt 0402_744765051A_5.1n 1 2
C1 1 N7 152.0253f
L1 1 N1 4.85n
L2 N1 N2 126.1185p
L3 N2 N3 129.1151p
L4 N3 N4 83.9388p
L5 N4 N5 48.3829p
L6 N5 N6 410.0049p
R1 2 N1 928.4837m
R2 2 N2 1.1544
R3 2 N3 936.8238m
R4 2 N4 762.4379m
R5 2 N5 638.6151m
R6 2 N6 365.9469m
R7 2 N7 1.9755
R8 2 1 1000000
.ends 0402_744765051A_5.1n
*******
.subckt 0402_744765051GA_5.1n 1 2
C1 1 N7 152.0253f
L1 1 N1 4.85n
L2 N1 N2 126.1185p
L3 N2 N3 129.1151p
L4 N3 N4 83.9388p
L5 N4 N5 48.3829p
L6 N5 N6 410.0049p
R1 2 N1 928.4837m
R2 2 N2 1.1544
R3 2 N3 936.8238m
R4 2 N4 762.4379m
R5 2 N5 638.6151m
R6 2 N6 365.9469m
R7 2 N7 1.9755
R8 2 1 1000000
.ends 0402_744765051GA_5.1n
*******
.subckt 0402_744765056A_5.6n 1 2
C1 1 N7 98.6102f
L1 1 N1 5.35n
L2 N1 N2 136.5935p
L3 N2 N3 134.3901p
L4 N3 N4 86.3994p
L5 N4 N5 49.4908p
L6 N5 N6 436.6862p
R1 2 N1 1.0593
R2 2 N2 1.2191
R3 2 N3 968.4352m
R4 2 N4 786.7350m
R5 2 N5 664.1795m
R6 2 N6 358.3856m
R7 2 N7 1.9734
R8 2 1 1000000
.ends 0402_744765056A_5.6n
*******
.subckt 0402_744765056GA_5.6n 1 2
C1 1 N7 98.6102f
L1 1 N1 5.35n
L2 N1 N2 136.5935p
L3 N2 N3 134.3901p
L4 N3 N4 86.3994p
L5 N4 N5 49.4908p
L6 N5 N6 436.6862p
R1 2 N1 1.0593
R2 2 N2 1.2191
R3 2 N3 968.4352m
R4 2 N4 786.7350m
R5 2 N5 664.1795m
R6 2 N6 358.3856m
R7 2 N7 1.9734
R8 2 1 1000000
.ends 0402_744765056GA_5.6n
*******
.subckt 0402_744765062A_6.2n 1 2
C1 1 N7 45.7108f
L1 1 N1 5.95n
L2 N1 N2 152.7755p
L3 N2 N3 145.7468p
L4 N3 N4 93.1160p
L5 N4 N5 52.7038p
L6 N5 N6 515.0878p
R1 2 N1 1.1816
R2 2 N2 1.3244
R3 2 N3 1.0501
R4 2 N4 860.9239m
R5 2 N5 743.2689m
R6 2 N6 348.3450m
R7 2 N7 1.9722
R8 2 1 1000000
.ends 0402_744765062A_6.2n
*******
.subckt 0402_744765062GA_6.2n 1 2
C1 1 N7 45.7108f
L1 1 N1 5.95n
L2 N1 N2 152.7755p
L3 N2 N3 145.7468p
L4 N3 N4 93.1160p
L5 N4 N5 52.7038p
L6 N5 N6 515.0878p
R1 2 N1 1.1816
R2 2 N2 1.3244
R3 2 N3 1.0501
R4 2 N4 860.9239m
R5 2 N5 743.2689m
R6 2 N6 348.3450m
R7 2 N7 1.9722
R8 2 1 1000000
.ends 0402_744765062GA_6.2n
*******
.subckt 0402_744765068A_6.8n 1 2
C1 1 N7 83.0836f
L1 1 N1 6.5n
L2 N1 N2 182.6013p
L3 N2 N3 191.0980p
L4 N3 N4 134.1514p
L5 N4 N5 72.1778p
L6 N5 N6 992.8975p
R1 2 N1 1.3834
R2 2 N2 1.7882
R3 2 N3 1.591
R4 2 N4 1.3965
R5 2 N5 1.3028
R6 2 N6 593.1976m
R7 2 N7 1.9678
R8 2 1 1000000
.ends 0402_744765068A_6.8n
*******
.subckt 0402_744765068GA_6.8n 1 2
C1 1 N7 83.0836f
L1 1 N1 6.5n
L2 N1 N2 182.6013p
L3 N2 N3 191.0980p
L4 N3 N4 134.1514p
L5 N4 N5 72.1778p
L6 N5 N6 992.8975p
R1 2 N1 1.3834
R2 2 N2 1.7882
R3 2 N3 1.591
R4 2 N4 1.3965
R5 2 N5 1.3028
R6 2 N6 593.1976m
R7 2 N7 1.9678
R8 2 1 1000000
.ends 0402_744765068GA_6.8n
*******
.subckt 0402_744765075A_7.5n 1 2
C1 1 N7 63.2462f
L1 1 N1 7.2n
L2 N1 N2 182.4916p
L3 N2 N3 191.0922p
L4 N3 N4 134.1543p
L5 N4 N5 72.1788p
L6 N5 N6 992.8935p
R1 2 N1 1.3798
R2 2 N2 1.7878
R3 2 N3 1.591
R4 2 N4 1.3965
R5 2 N5 1.3028
R6 2 N6 592.9804m
R7 2 N7 1.9677
R8 2 1 1000000
.ends 0402_744765075A_7.5n
*******
.subckt 0402_744765075GA_7.5n 1 2
C1 1 N7 63.2462f
L1 1 N1 7.2n
L2 N1 N2 182.4916p
L3 N2 N3 191.0922p
L4 N3 N4 134.1543p
L5 N4 N5 72.1788p
L6 N5 N6 992.8935p
R1 2 N1 1.3798
R2 2 N2 1.7878
R3 2 N3 1.591
R4 2 N4 1.3965
R5 2 N5 1.3028
R6 2 N6 592.9804m
R7 2 N7 1.9677
R8 2 1 1000000
.ends 0402_744765075GA_7.5n
*******
.subckt 0402_744765082A_8.2n 1 2
C1 1 N7 78.4949f
L1 1 N1 7.8n
L2 N1 N2 182.4916p
L3 N2 N3 191.0922p
L4 N3 N4 135.1153p
L5 N4 N5 72.4800p
L6 N5 N6 992.8935p
R1 2 N1 1.5865
R2 2 N2 1.8494
R3 2 N3 1.6039
R4 2 N4 1.4003
R5 2 N5 1.3046
R6 2 N6 570.0508m
R7 2 N7 1.9656
R8 2 1 1000000
.ends 0402_744765082A_8.2n
*******
.subckt 0402_744765082GA_8.2n 1 2
C1 1 N7 78.4949f
L1 1 N1 7.8n
L2 N1 N2 182.4916p
L3 N2 N3 191.0922p
L4 N3 N4 135.1153p
L5 N4 N5 72.4800p
L6 N5 N6 992.8935p
R1 2 N1 1.5865
R2 2 N2 1.8494
R3 2 N3 1.6039
R4 2 N4 1.4003
R5 2 N5 1.3046
R6 2 N6 570.0508m
R7 2 N7 1.9656
R8 2 1 1000000
.ends 0402_744765082GA_8.2n
*******
.subckt 0402_744765087A_8.7n 1 2
C1 1 N7 22.0581f
L1 1 N1 8.3n
L2 N1 N2 155.0829p
L3 N2 N3 183.5830p
L4 N3 N4 207.6467p
L5 N4 N5 101.7920p
L6 N5 N6 992.8935p
R1 2 N1 3.3489
R2 2 N2 2.9363
R3 2 N3 2.4492
R4 2 N4 2.0775
R5 2 N5 1.9055
R6 2 N6 644.9946m
R7 2 N7 1.9366
R8 2 1 1000000
.ends 0402_744765087A_8.7n
*******
.subckt 0402_744765090A_9n 1 2
C1 1 N7 49.9561f
L1 1 N1 8.55n
L2 N1 N2 94.0460p
L3 N2 N3 158.0317p
L4 N3 N4 203.1479p
L5 N4 N5 100.8256p
L6 N5 N6 976.1723p
R1 2 N1 3.1128
R2 2 N2 2.6843
R3 2 N3 2.3587
R4 2 N4 2.0602
R5 2 N5 1.894
R6 2 N6 619.8332m
R7 2 N7 1.9341
R8 2 1 1000000
.ends 0402_744765090A_9n
*******
.subckt 0402_744765090GA_9n 1 2
C1 1 N7 49.9561f
L1 1 N1 8.55n
L2 N1 N2 94.0460p
L3 N2 N3 158.0317p
L4 N3 N4 203.1479p
L5 N4 N5 100.8256p
L6 N5 N6 976.1723p
R1 2 N1 3.1128
R2 2 N2 2.6843
R3 2 N3 2.3587
R4 2 N4 2.0602
R5 2 N5 1.894
R6 2 N6 619.8332m
R7 2 N7 1.9341
R8 2 1 1000000
.ends 0402_744765090GA_9n
*******
.subckt 0402_744765095A_9.5n 1 2
C1 1 N7 22.0867f
L1 1 N1 9n
L2 N1 N2 140.7895p
L3 N2 N3 192.8702p
L4 N3 N4 213.0035p
L5 N4 N5 165.7744p
L6 N5 N6 1.0059n
R1 2 N1 2.9812
R2 2 N2 3.6414
R3 2 N3 3.7736
R4 2 N4 3.2115
R5 2 N5 2.8792
R6 2 N6 1.1524
R7 2 N7 1.9144
R8 2 1 1000000
.ends 0402_744765095A_9.5n
*******
.subckt 0402_744765095GA_9.5n 1 2
C1 1 N7 22.0867f
L1 1 N1 9n
L2 N1 N2 140.7895p
L3 N2 N3 192.8702p
L4 N3 N4 213.0035p
L5 N4 N5 165.7744p
L6 N5 N6 1.0059n
R1 2 N1 2.9812
R2 2 N2 3.6414
R3 2 N3 3.7736
R4 2 N4 3.2115
R5 2 N5 2.8792
R6 2 N6 1.1524
R7 2 N7 1.9144
R8 2 1 1000000
.ends 0402_744765095GA_9.5n
*******
.subckt 0402_744765110A_10n 1 2
C1 1 N7 21.8477f
L1 1 N1 9.5n
L2 N1 N2 93.1599p
L3 N2 N3 111.5855p
L4 N3 N4 164.2473p
L5 N4 N5 175.9956p
L6 N5 N6 315.8247p
R1 2 N1 3.0555
R2 2 N2 4.1558
R3 2 N3 4.0385
R4 2 N4 3.3362
R5 2 N5 2.8717
R6 2 N6 1.0146
R7 2 N7 4.69
R8 2 1 1000000
.ends 0402_744765110A_10n
*******
.subckt 0402_744765110GA_10n 1 2
C1 1 N7 21.8477f
L1 1 N1 9.5n
L2 N1 N2 93.1599p
L3 N2 N3 111.5855p
L4 N3 N4 164.2473p
L5 N4 N5 175.9956p
L6 N5 N6 315.8247p
R1 2 N1 3.0555
R2 2 N2 4.1558
R3 2 N3 4.0385
R4 2 N4 3.3362
R5 2 N5 2.8717
R6 2 N6 1.0146
R7 2 N7 4.69
R8 2 1 1000000
.ends 0402_744765110GA_10n
*******
.subckt 0402_744765111A_11n 1 2
C1 1 N7 103.8026f
L1 1 N1 10.5n
L2 N1 N2 107.8041p
L3 N2 N3 139.0629p
L4 N3 N4 187.4208p
L5 N4 N5 187.7668p
L6 N5 N6 562.0267p
R1 2 N1 2.5853
R2 2 N2 3.8634
R3 2 N3 3.787
R4 2 N4 3.0854
R5 2 N5 2.6663
R6 2 N6 679.0439m
R7 2 N7 3.6956
R8 2 1 1000000
.ends 0402_744765111A_11n
*******
.subckt 0402_744765111GA_11n 1 2
C1 1 N7 103.8026f
L1 1 N1 10.5n
L2 N1 N2 107.8041p
L3 N2 N3 139.0629p
L4 N3 N4 187.4208p
L5 N4 N5 187.7668p
L6 N5 N6 562.0267p
R1 2 N1 2.5853
R2 2 N2 3.8634
R3 2 N3 3.787
R4 2 N4 3.0854
R5 2 N5 2.6663
R6 2 N6 679.0439m
R7 2 N7 3.6956
R8 2 1 1000000
.ends 0402_744765111GA_11n
*******
.subckt 0402_744765112A_12n 1 2
C1 1 N7 96.6372f
L1 1 N1 11.4n
L2 N1 N2 143.4175p
L3 N2 N3 164.4827p
L4 N3 N4 198.3812p
L5 N4 N5 190.1172p
L6 N5 N6 566.2931p
R1 2 N1 2.8587
R2 2 N2 3.9879
R3 2 N3 3.8628
R4 2 N4 3.1168
R5 2 N5 2.6705
R6 2 N6 620.5290m
R7 2 N7 3.6931
R8 2 1 1000000
.ends 0402_744765112A_12n
*******
.subckt 0402_744765112GA_12n 1 2
C1 1 N7 96.6372f
L1 1 N1 11.4n
L2 N1 N2 143.4175p
L3 N2 N3 164.4827p
L4 N3 N4 198.3812p
L5 N4 N5 190.1172p
L6 N5 N6 566.2931p
R1 2 N1 2.8587
R2 2 N2 3.9879
R3 2 N3 3.8628
R4 2 N4 3.1168
R5 2 N5 2.6705
R6 2 N6 620.5290m
R7 2 N7 3.6931
R8 2 1 1000000
.ends 0402_744765112GA_12n
*******
.subckt 0402_744765113A_13n 1 2
C1 1 N7 100.7608f
L1 1 N1 12.4n
L2 N1 N2 178.9608p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 195.4094p
L6 N5 N6 746.9179p
R1 2 N1 3.1102
R2 2 N2 4.1255
R3 2 N3 3.9536
R4 2 N4 3.1755
R5 2 N5 2.7066
R6 2 N6 715.2736m
R7 2 N7 3.6906
R8 2 1 1000000
.ends 0402_744765113A_13n
*******
.subckt 0402_744765113GA_13n 1 2
C1 1 N7 100.7608f
L1 1 N1 12.4n
L2 N1 N2 178.9608p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 195.4094p
L6 N5 N6 746.9179p
R1 2 N1 3.1102
R2 2 N2 4.1255
R3 2 N3 3.9536
R4 2 N4 3.1755
R5 2 N5 2.7066
R6 2 N6 715.2736m
R7 2 N7 3.6906
R8 2 1 1000000
.ends 0402_744765113GA_13n
*******
.subckt 0402_744765115A_15n 1 2
C1 1 N7 78.1968f
L1 1 N1 14.3n
L2 N1 N2 184.4580p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 206.5524p
L6 N5 N6 986.2845p
R1 2 N1 3.7539
R2 2 N2 4.5237
R3 2 N3 4.1991
R4 2 N4 3.3195
R5 2 N5 2.7862
R6 2 N6 695.4261m
R7 2 N7 3.6817
R8 2 1 1000000
.ends 0402_744765115A_15n
*******
.subckt 0402_744765115GA_15n 1 2
C1 1 N7 78.1968f
L1 1 N1 14.3n
L2 N1 N2 184.4580p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 206.5524p
L6 N5 N6 986.2845p
R1 2 N1 3.7539
R2 2 N2 4.5237
R3 2 N3 4.1991
R4 2 N4 3.3195
R5 2 N5 2.7862
R6 2 N6 695.4261m
R7 2 N7 3.6817
R8 2 1 1000000
.ends 0402_744765115GA_15n
*******
.subckt 0402_744765116A_16n 1 2
C1 1 N7 89.6533f
L1 1 N1 15.2n
L2 N1 N2 184.4580p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 206.5663p
L6 N5 N6 986.1019p
R1 2 N1 3.7549
R2 2 N2 4.5245
R3 2 N3 4.1995
R4 2 N4 3.3196
R5 2 N5 2.7862
R6 2 N6 694.1841m
R7 2 N7 3.6818
R8 2 1 1000000
.ends 0402_744765116A_16n
*******
.subckt 0402_744765116GA_16n 1 2
C1 1 N7 89.6533f
L1 1 N1 15.2n
L2 N1 N2 184.4580p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 206.5663p
L6 N5 N6 986.1019p
R1 2 N1 3.7549
R2 2 N2 4.5245
R3 2 N3 4.1995
R4 2 N4 3.3196
R5 2 N5 2.7862
R6 2 N6 694.1841m
R7 2 N7 3.6818
R8 2 1 1000000
.ends 0402_744765116GA_16n
*******
.subckt 0402_744765118A_18n 1 2
C1 1 N7 82.8466f
L1 1 N1 17.3n
L2 N1 N2 184.4580p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 209.5938p
L6 N5 N6 863.2763p
R1 2 N1 4.0095
R2 2 N2 4.7252
R3 2 N3 4.2808
R4 2 N4 3.3605
R5 2 N5 2.7684
R6 2 N6 265.8437m
R7 2 N7 3.677
R8 2 1 1000000
.ends 0402_744765118A_18n
*******
.subckt 0402_744765118GA_18n 1 2
C1 1 N7 82.8466f
L1 1 N1 17.3n
L2 N1 N2 184.4580p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 209.5938p
L6 N5 N6 863.2763p
R1 2 N1 4.0095
R2 2 N2 4.7252
R3 2 N3 4.2808
R4 2 N4 3.3605
R5 2 N5 2.7684
R6 2 N6 265.8437m
R7 2 N7 3.677
R8 2 1 1000000
.ends 0402_744765118GA_18n
*******
.subckt 0402_744765119A_19n 1 2
C1 1 N7 71.0935f
L1 1 N1 18n
L2 N1 N2 184.4421p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 261.9862p
L6 N5 N6 994.6071p
R1 2 N1 7.3531
R2 2 N2 8.1557
R3 2 N3 4.2808
R4 2 N4 3.6212
R5 2 N5 2.9318
R6 2 N6 1.1848
R7 2 N7 3.6102
R8 2 1 1000000
.ends 0402_744765119A_19n
*******
.subckt 0402_744765119GA_19n 1 2
C1 1 N7 71.0935f
L1 1 N1 18n
L2 N1 N2 184.4421p
L3 N2 N3 191.2043p
L4 N3 N4 212.1927p
L5 N4 N5 261.9862p
L6 N5 N6 994.6071p
R1 2 N1 7.3531
R2 2 N2 8.1557
R3 2 N3 4.2808
R4 2 N4 3.6212
R5 2 N5 2.9318
R6 2 N6 1.1848
R7 2 N7 3.6102
R8 2 1 1000000
.ends 0402_744765119GA_19n
*******
.subckt 0402_744765120A_20n 1 2
C1 1 N7 82.0086f
L1 1 N1 19.2n
L2 N1 N2 351.8529p
L3 N2 N3 569.0964p
L4 N3 N4 651.0460p
L5 N4 N5 573.2864p
L6 N5 N6 1.1149n
R1 2 N1 3.9611
R2 2 N2 4.7233
R3 2 N3 4.3048
R4 2 N4 3.4051
R5 2 N5 2.8219
R6 2 N6 856.8275m
R7 2 N7 3.6791
R8 2 1 1000000
.ends 0402_744765120A_20n
*******
.subckt 0402_744765120GA_20n 1 2
C1 1 N7 82.0086f
L1 1 N1 19.2n
L2 N1 N2 351.8529p
L3 N2 N3 569.0964p
L4 N3 N4 651.0460p
L5 N4 N5 573.2864p
L6 N5 N6 1.1149n
R1 2 N1 3.9611
R2 2 N2 4.7233
R3 2 N3 4.3048
R4 2 N4 3.4051
R5 2 N5 2.8219
R6 2 N6 856.8275m
R7 2 N7 3.6791
R8 2 1 1000000
.ends 0402_744765120GA_20n
*******
.subckt 0402_744765122A_22n 1 2
C1 1 N7 69.0722f
L1 1 N1 21.2n
L2 N1 N2 432.7651p
L3 N2 N3 416.8593p
L4 N3 N4 516.5121p
L5 N4 N5 519.8417p
L6 N5 N6 1.1021n
R1 2 N1 3.9788
R2 2 N2 4.7174
R3 2 N3 4.2842
R4 2 N4 3.3872
R5 2 N5 2.809
R6 2 N6 789.1994m
R7 2 N7 3.6755
R8 2 1 1000000
.ends 0402_744765122A_22n
*******
.subckt 0402_744765122GA_22n 1 2
C1 1 N7 69.0722f
L1 1 N1 21.2n
L2 N1 N2 432.7651p
L3 N2 N3 416.8593p
L4 N3 N4 516.5121p
L5 N4 N5 519.8417p
L6 N5 N6 1.1021n
R1 2 N1 3.9788
R2 2 N2 4.7174
R3 2 N3 4.2842
R4 2 N4 3.3872
R5 2 N5 2.809
R6 2 N6 789.1994m
R7 2 N7 3.6755
R8 2 1 1000000
.ends 0402_744765122GA_22n
*******
.subckt 0402_744765123A_23n 1 2
C1 1 N7 76.1232f
L1 1 N1 22.2n
L2 N1 N2 603.2051p
L3 N2 N3 463.5833p
L4 N3 N4 525.9776p
L5 N4 N5 526.0674p
L6 N5 N6 1.1066n
R1 2 N1 4.0071
R2 2 N2 4.7258
R3 2 N3 4.2862
R4 2 N4 3.3881
R5 2 N5 2.8101
R6 2 N6 791.9371m
R7 2 N7 3.6775
R8 2 1 1000000
.ends 0402_744765123A_23n
*******
.subckt 0402_744765123GA_23n 1 2
C1 1 N7 76.1232f
L1 1 N1 22.2n
L2 N1 N2 603.2051p
L3 N2 N3 463.5833p
L4 N3 N4 525.9776p
L5 N4 N5 526.0674p
L6 N5 N6 1.1066n
R1 2 N1 4.0071
R2 2 N2 4.7258
R3 2 N3 4.2862
R4 2 N4 3.3881
R5 2 N5 2.8101
R6 2 N6 791.9371m
R7 2 N7 3.6775
R8 2 1 1000000
.ends 0402_744765123GA_23n
*******
.subckt 0402_744765124A_24n 1 2
C1 1 N7 80.2086f
L1 1 N1 23.2n
L2 N1 N2 599.8434p
L3 N2 N3 663.0589p
L4 N3 N4 866.2427p
L5 N4 N5 801.8895p
L6 N5 N6 1.2620n
R1 2 N1 3.9944
R2 2 N2 4.7297
R3 2 N3 4.3203
R4 2 N4 3.4491
R5 2 N5 2.8737
R6 2 N6 1.0405
R7 2 N7 3.6857
R8 2 1 1000000
.ends 0402_744765124A_24n
*******
.subckt 0402_744765124GA_24n 1 2
C1 1 N7 80.2086f
L1 1 N1 23.2n
L2 N1 N2 599.8434p
L3 N2 N3 663.0589p
L4 N3 N4 866.2427p
L5 N4 N5 801.8895p
L6 N5 N6 1.2620n
R1 2 N1 3.9944
R2 2 N2 4.7297
R3 2 N3 4.3203
R4 2 N4 3.4491
R5 2 N5 2.8737
R6 2 N6 1.0405
R7 2 N7 3.6857
R8 2 1 1000000
.ends 0402_744765124GA_24n
*******
.subckt 0402_744765127A_27n 1 2
C1 1 N7 70.9595f
L1 1 N1 26n
L2 N1 N2 731.7231p
L3 N2 N3 692.2963p
L4 N3 N4 867.5511p
L5 N4 N5 803.8989p
L6 N5 N6 1.2638n
R1 2 N1 4.0219
R2 2 N2 4.7397
R3 2 N3 4.3216
R4 2 N4 3.4494
R5 2 N5 2.8743
R6 2 N6 1.042
R7 2 N7 3.6834
R8 2 1 1000000
.ends 0402_744765127A_27n
*******
.subckt 0402_744765127GA_27n 1 2
C1 1 N7 70.9595f
L1 1 N1 26n
L2 N1 N2 731.7231p
L3 N2 N3 692.2963p
L4 N3 N4 867.5511p
L5 N4 N5 803.8989p
L6 N5 N6 1.2638n
R1 2 N1 4.0219
R2 2 N2 4.7397
R3 2 N3 4.3216
R4 2 N4 3.4494
R5 2 N5 2.8743
R6 2 N6 1.042
R7 2 N7 3.6834
R8 2 1 1000000
.ends 0402_744765127GA_27n
*******
.subckt 0402_744765130A_30n 1 2
C1 1 N7 74.1373f
L1 1 N1 29.1n
L2 N1 N2 1.1419n
L3 N2 N3 791.8263p
L4 N3 N4 1.3275n
L5 N4 N5 1.1844n
L6 N5 N6 1.4598n
R1 2 N1 4.7216
R2 2 N2 4.7246
R3 2 N3 4.3857
R4 2 N4 3.5901
R5 2 N5 3.02
R6 2 N6 1.5055
R7 2 N7 3.7342
R8 2 1 1000000
.ends 0402_744765130A_30n
*******
.subckt 0402_744765130GA_30n 1 2
C1 1 N7 74.1373f
L1 1 N1 29.1n
L2 N1 N2 1.1419n
L3 N2 N3 791.8263p
L4 N3 N4 1.3275n
L5 N4 N5 1.1844n
L6 N5 N6 1.4598n
R1 2 N1 4.7216
R2 2 N2 4.7246
R3 2 N3 4.3857
R4 2 N4 3.5901
R5 2 N5 3.02
R6 2 N6 1.5055
R7 2 N7 3.7342
R8 2 1 1000000
.ends 0402_744765130GA_30n
*******
.subckt 0402_744765133A_33n 1 2
C1 1 N7 64.5625f
L1 1 N1 32.2n
L2 N1 N2 1.0670n
L3 N2 N3 301.7329p
L4 N3 N4 1.1241n
L5 N4 N5 1.1159n
L6 N5 N6 1.4412n
R1 2 N1 4.9858
R2 2 N2 4.6172
R3 2 N3 4.2824
R4 2 N4 3.5281
R5 2 N5 2.9667
R6 2 N6 1.3303
R7 2 N7 3.7565
R8 2 1 1000000
.ends 0402_744765133A_33n
*******
.subckt 0402_744765133GA_33n 1 2
C1 1 N7 64.5625f
L1 1 N1 32.2n
L2 N1 N2 1.0670n
L3 N2 N3 301.7329p
L4 N3 N4 1.1241n
L5 N4 N5 1.1159n
L6 N5 N6 1.4412n
R1 2 N1 4.9858
R2 2 N2 4.6172
R3 2 N3 4.2824
R4 2 N4 3.5281
R5 2 N5 2.9667
R6 2 N6 1.3303
R7 2 N7 3.7565
R8 2 1 1000000
.ends 0402_744765133GA_33n
*******
.subckt 0402_744765136A_36n 1 2
C1 1 N7 66.7653f
L1 1 N1 35n
L2 N1 N2 1.5270n
L3 N2 N3 575.4741p
L4 N3 N4 1.2818n
L5 N4 N5 1.1948n
L6 N5 N6 1.4721n
R1 2 N1 5.0899
R2 2 N2 4.6682
R3 2 N3 4.3299
R4 2 N4 3.5641
R5 2 N5 2.9915
R6 2 N6 1.3748
R7 2 N7 3.7626
R8 2 1 1000000
.ends 0402_744765136A_36n
*******
.subckt 0402_744765136GA_36n 1 2
C1 1 N7 66.7653f
L1 1 N1 35n
L2 N1 N2 1.5270n
L3 N2 N3 575.4741p
L4 N3 N4 1.2818n
L5 N4 N5 1.1948n
L6 N5 N6 1.4721n
R1 2 N1 5.0899
R2 2 N2 4.6682
R3 2 N3 4.3299
R4 2 N4 3.5641
R5 2 N5 2.9915
R6 2 N6 1.3748
R7 2 N7 3.7626
R8 2 1 1000000
.ends 0402_744765136GA_36n
*******
.subckt 0402_744765139A_39n 1 2
C1 1 N7 57.6983f
L1 1 N1 37n
L2 N1 N2 1.3611n
L3 N2 N3 1.7441n
L4 N3 N4 2.0947n
L5 N4 N5 2.0539n
L6 N5 N6 1.8246n
R1 2 N1 6.5863
R2 2 N2 4.7459
R3 2 N3 4.782
R4 2 N4 4.0992
R5 2 N5 3.4699
R6 2 N6 2.3704
R7 2 N7 3.9032
R8 2 1 1000000
.ends 0402_744765139A_39n
*******
.subckt 0402_744765139GA_39n 1 2
C1 1 N7 57.6983f
L1 1 N1 37n
L2 N1 N2 1.3611n
L3 N2 N3 1.7441n
L4 N3 N4 2.0947n
L5 N4 N5 2.0539n
L6 N5 N6 1.8246n
R1 2 N1 6.5863
R2 2 N2 4.7459
R3 2 N3 4.782
R4 2 N4 4.0992
R5 2 N5 3.4699
R6 2 N6 2.3704
R7 2 N7 3.9032
R8 2 1 1000000
.ends 0402_744765139GA_39n
*******
.subckt 0402_744765140A_40n 1 2
C1 1 N7 66.0474f
L1 1 N1 38n
L2 N1 N2 1.3721n
L3 N2 N3 1.7430n
L4 N3 N4 2.0947n
L5 N4 N5 2.0540n
L6 N5 N6 1.8246n
R1 2 N1 6.5922
R2 2 N2 4.7457
R3 2 N3 4.7819
R4 2 N4 4.0993
R5 2 N5 3.47
R6 2 N6 2.3705
R7 2 N7 3.9045
R8 2 1 1000000
.ends 0402_744765140A_40n
*******
.subckt 0402_744765140GA_40n 1 2
C1 1 N7 66.0474f
L1 1 N1 38n
L2 N1 N2 1.3721n
L3 N2 N3 1.7430n
L4 N3 N4 2.0947n
L5 N4 N5 2.0540n
L6 N5 N6 1.8246n
R1 2 N1 6.5922
R2 2 N2 4.7457
R3 2 N3 4.7819
R4 2 N4 4.0993
R5 2 N5 3.47
R6 2 N6 2.3705
R7 2 N7 3.9045
R8 2 1 1000000
.ends 0402_744765140GA_40n
*******
.subckt 0402_744765143A_43n 1 2
C1 1 N7 63.9382f
L1 1 N1 40n
L2 N1 N2 1.4956n
L3 N2 N3 344.8851p
L4 N3 N4 1.5260n
L5 N4 N5 1.7872n
L6 N5 N6 1.7511n
R1 2 N1 7.011
R2 2 N2 4.1838
R3 2 N3 4.3654
R4 2 N4 3.8612
R5 2 N5 3.3237
R6 2 N6 2.1834
R7 2 N7 3.9867
R8 2 1 1000000
.ends 0402_744765143A_43n
*******
.subckt 0402_744765143GA_43n 1 2
C1 1 N7 63.9382f
L1 1 N1 40n
L2 N1 N2 1.4956n
L3 N2 N3 344.8851p
L4 N3 N4 1.5260n
L5 N4 N5 1.7872n
L6 N5 N6 1.7511n
R1 2 N1 7.011
R2 2 N2 4.1838
R3 2 N3 4.3654
R4 2 N4 3.8612
R5 2 N5 3.3237
R6 2 N6 2.1834
R7 2 N7 3.9867
R8 2 1 1000000
.ends 0402_744765143GA_43n
*******
.subckt 0402_744765147A_47n 1 2
C1 1 N7 0.122209180174463p
L1 1 N1 47n
L2 N1 N2 1.7547n
L3 N2 N3 1.8894n
L4 N3 N4 1.9412n
L5 N4 N5 1.2813n
L6 N5 N6 1.3683n
R1 2 N1 7.3009
R2 2 N2 4.7788
R3 2 N3 4.5418
R4 2 N4 3.7494
R5 2 N5 3.1902
R6 2 N6 2.1172
R7 2 N7 4.0266
R8 2 1 1000000
.ends 0402_744765147A_47n
*******
.subckt 0402_744765147GA_47n 1 2
C1 1 N7 0.122209180174463p
L1 1 N1 47n
L2 N1 N2 1.7547n
L3 N2 N3 1.8894n
L4 N3 N4 1.9412n
L5 N4 N5 1.2813n
L6 N5 N6 1.3683n
R1 2 N1 7.3009
R2 2 N2 4.7788
R3 2 N3 4.5418
R4 2 N4 3.7494
R5 2 N5 3.1902
R6 2 N6 2.1172
R7 2 N7 4.0266
R8 2 1 1000000
.ends 0402_744765147GA_47n
*******
.subckt 0402_744765151A_51n 1 2
C1 1 N7 0.162178770866817p
L1 1 N1 49n
L2 N1 N2 1.8328n
L3 N2 N3 1.8613n
L4 N3 N4 2.0899n
L5 N4 N5 1.4179n
L6 N5 N6 1.4248n
R1 2 N1 8.9988
R2 2 N2 4.9103
R3 2 N3 4.5655
R4 2 N4 3.85
R5 2 N5 3.3016
R6 2 N6 2.3014
R7 2 N7 4.2769
R8 2 1 1000000
.ends 0402_744765151A_51n
*******
.subckt 0402_744765151GA_51n 1 2
C1 1 N7 0.162178770866817p
L1 1 N1 49n
L2 N1 N2 1.8328n
L3 N2 N3 1.8613n
L4 N3 N4 2.0899n
L5 N4 N5 1.4179n
L6 N5 N6 1.4248n
R1 2 N1 8.9988
R2 2 N2 4.9103
R3 2 N3 4.5655
R4 2 N4 3.85
R5 2 N5 3.3016
R6 2 N6 2.3014
R7 2 N7 4.2769
R8 2 1 1000000
.ends 0402_744765151GA_51n
*******
.subckt 0402_744765156A_56n 1 2
C1 1 N7 0.146024899315836p
L1 1 N1 56n
L2 N1 N2 1.8359n
L3 N2 N3 1.9056n
L4 N3 N4 2.0899n
L5 N4 N5 1.6907n
L6 N5 N6 1.5178n
R1 2 N1 10.2892
R2 2 N2 5.7153
R3 2 N3 4.8061
R4 2 N4 4.0222
R5 2 N5 3.4372
R6 2 N6 2.464
R7 2 N7 4.5128
R8 2 1 1000000
.ends 0402_744765156A_56n
*******
.subckt 0402_744765156GA_56n 1 2
C1 1 N7 0.146024899315836p
L1 1 N1 56n
L2 N1 N2 1.8359n
L3 N2 N3 1.9056n
L4 N3 N4 2.0899n
L5 N4 N5 1.6907n
L6 N5 N6 1.5178n
R1 2 N1 10.2892
R2 2 N2 5.7153
R3 2 N3 4.8061
R4 2 N4 4.0222
R5 2 N5 3.4372
R6 2 N6 2.464
R7 2 N7 4.5128
R8 2 1 1000000
.ends 0402_744765156GA_56n
*******
.subckt 0402_744765168A_68n 1 2
C1 1 N7 0.14193886767822p
L1 1 N1 68n
L2 N1 N2 1.8359n
L3 N2 N3 1.9051n
L4 N3 N4 2.0899n
L5 N4 N5 2.0603n
L6 N5 N6 1.8507n
R1 2 N1 14.1035
R2 2 N2 10.1194
R3 2 N3 6.2545
R4 2 N4 4.8005
R5 2 N5 3.9377
R6 2 N6 2.6435
R7 2 N7 5.4165
R8 2 1 1000000
.ends 0402_744765168A_68n
*******
.subckt 0402_744765168GA_68n 1 2
C1 1 N7 0.14193886767822p
L1 1 N1 68n
L2 N1 N2 1.8359n
L3 N2 N3 1.9051n
L4 N3 N4 2.0899n
L5 N4 N5 2.0603n
L6 N5 N6 1.8507n
R1 2 N1 14.1035
R2 2 N2 10.1194
R3 2 N3 6.2545
R4 2 N4 4.8005
R5 2 N5 3.9377
R6 2 N6 2.6435
R7 2 N7 5.4165
R8 2 1 1000000
.ends 0402_744765168GA_68n
*******
.subckt 0402_744765175A_75n 1 2
C1 1 N7 0.14057743614158p
L1 1 N1 73n
L2 N1 N2 2.1879n
L3 N2 N3 1.9195n
L4 N3 N4 3.2201n
L5 N4 N5 2.9613n
L6 N5 N6 2.2215n
R1 2 N1 14.3027
R2 2 N2 10.0124
R3 2 N3 6.2565
R4 2 N4 4.806
R5 2 N5 3.9428
R6 2 N6 2.6498
R7 2 N7 5.4161
R8 2 1 1000000
.ends 0402_744765175A_75n
*******
.subckt 0402_744765175GA_75n 1 2
C1 1 N7 0.14057743614158p
L1 1 N1 73n
L2 N1 N2 2.1879n
L3 N2 N3 1.9195n
L4 N3 N4 3.2201n
L5 N4 N5 2.9613n
L6 N5 N6 2.2215n
R1 2 N1 14.3027
R2 2 N2 10.0124
R3 2 N3 6.2565
R4 2 N4 4.806
R5 2 N5 3.9428
R6 2 N6 2.6498
R7 2 N7 5.4161
R8 2 1 1000000
.ends 0402_744765175GA_75n
*******
.subckt 0402_744765182A_82n 1 2
C1 1 N7 0.137291581435019p
L1 1 N1 77n
L2 N1 N2 2.3273n
L3 N2 N3 1.7144n
L4 N3 N4 5.3645n
L5 N4 N5 4.1000n
L6 N5 N6 2.6484n
R1 2 N1 16.6704
R2 2 N2 10.1574
R3 2 N3 6.2692
R4 2 N4 4.8192
R5 2 N5 3.9544
R6 2 N6 2.668
R7 2 N7 5.4281
R8 2 1 1000000
.ends 0402_744765182A_82n
*******
.subckt 0402_744765182GA_82n 1 2
C1 1 N7 0.137291581435019p
L1 1 N1 77n
L2 N1 N2 2.3273n
L3 N2 N3 1.7144n
L4 N3 N4 5.3645n
L5 N4 N5 4.1000n
L6 N5 N6 2.6484n
R1 2 N1 16.6704
R2 2 N2 10.1574
R3 2 N3 6.2692
R4 2 N4 4.8192
R5 2 N5 3.9544
R6 2 N6 2.668
R7 2 N7 5.4281
R8 2 1 1000000
.ends 0402_744765182GA_82n
*******
.subckt 0402_744765191A_91n 1 2
C1 1 N7 0.152732460692871p
L1 1 N1 84n
L2 N1 N2 2.4371n
L3 N2 N3 2.7767n
L4 N3 N4 6.3842n
L5 N4 N5 4.9583n
L6 N5 N6 2.9884n
R1 2 N1 16.6013
R2 2 N2 10.3446
R3 2 N3 6.2755
R4 2 N4 4.831
R5 2 N5 3.9671
R6 2 N6 2.6894
R7 2 N7 5.4287
R8 2 1 1000000
.ends 0402_744765191A_91n
*******
.subckt 0402_744765191GA_91n 1 2
C1 1 N7 0.152732460692871p
L1 1 N1 84n
L2 N1 N2 2.4371n
L3 N2 N3 2.7767n
L4 N3 N4 6.3842n
L5 N4 N5 4.9583n
L6 N5 N6 2.9884n
R1 2 N1 16.6013
R2 2 N2 10.3446
R3 2 N3 6.2755
R4 2 N4 4.831
R5 2 N5 3.9671
R6 2 N6 2.6894
R7 2 N7 5.4287
R8 2 1 1000000
.ends 0402_744765191GA_91n
*******
.subckt 0402_744765210A_100n 1 2
C1 1 N7 0.149883412868408p
L1 1 N1 90n
L2 N1 N2 2.4584n
L3 N2 N3 2.8416n
L4 N3 N4 6.4448n
L5 N4 N5 5.0217n
L6 N5 N6 3.0148n
R1 2 N1 16.5885
R2 2 N2 10.3651
R3 2 N3 6.2758
R4 2 N4 4.832
R5 2 N5 3.9682
R6 2 N6 2.6912
R7 2 N7 5.4285
R8 2 1 1000000
.ends 0402_744765210A_100n
*******
.subckt 0402_744765210GA_100n 1 2
C1 1 N7 0.149883412868408p
L1 1 N1 90n
L2 N1 N2 2.4584n
L3 N2 N3 2.8416n
L4 N3 N4 6.4448n
L5 N4 N5 5.0217n
L6 N5 N6 3.0148n
R1 2 N1 16.5885
R2 2 N2 10.3651
R3 2 N3 6.2758
R4 2 N4 4.832
R5 2 N5 3.9682
R6 2 N6 2.6912
R7 2 N7 5.4285
R8 2 1 1000000
.ends 0402_744765210GA_100n
*******
.subckt 0402_744765212A_120n 1 2
C1 1 N7 0.174451079715985p
L1 1 N1 108n
L2 N1 N2 4.1236n
L3 N2 N3 3.8718n
L4 N3 N4 10.5290n
L5 N4 N5 7.8997n
L6 N5 N6 4.0651n
R1 2 N1 17.611
R2 2 N2 10.2045
R3 2 N3 6.2999
R4 2 N4 4.8859
R5 2 N5 4.0186
R6 2 N6 2.7737
R7 2 N7 5.4338
R8 2 1 1000000
.ends 0402_744765212A_120n
*******
.subckt 0402_744765212GA_120n 1 2
C1 1 N7 0.174451079715985p
L1 1 N1 108n
L2 N1 N2 4.1236n
L3 N2 N3 3.8718n
L4 N3 N4 10.5290n
L5 N4 N5 7.8997n
L6 N5 N6 4.0651n
R1 2 N1 17.611
R2 2 N2 10.2045
R3 2 N3 6.2999
R4 2 N4 4.8859
R5 2 N5 4.0186
R6 2 N6 2.7737
R7 2 N7 5.4338
R8 2 1 1000000
.ends 0402_744765212GA_120n
*******
.subckt 0603_744761016A_1.6n 1 2
C1 1 N7 0.101321187099044p
L1 1 N1 1.5n
L2 N1 N2 46.4315p
L3 N2 N3 24.9647p
L4 N3 N4 99.4232p
L5 N4 N5 75.1462p
L6 N5 N6 53.5367p
R1 2 N1 364.8342m
R2 2 N2 426.2027m
R3 2 N3 95.2027m
R4 2 N4 110.1936m
R5 2 N5 95.0487m
R6 2 N6 87.4456m
R7 2 N7 1.946
R8 2 1 1000000
.ends 0603_744761016A_1.6n
*******
.subckt 0603_744761018A_1.8n 1 2
C1 1 N7 0.0900632774213724p
L1 1 N1 1.7n
L2 N1 N2 86.9703p
L3 N2 N3 70.3590p
L4 N3 N4 138.1753p
L5 N4 N5 75.3428p
L6 N5 N6 53.5940p
R1 2 N1 438.5420m
R2 2 N2 420.7053m
R3 2 N3 141.6519m
R4 2 N4 133.7273m
R5 2 N5 113.6405m
R6 2 N6 87.6297m
R7 2 N7 1.946
R8 2 1 1000000
.ends 0603_744761018A_1.8n
*******
.subckt 0603_744761020A_2n 1 2
C1 1 N7 0.26601865968033p
L1 1 N1 1.8n
L2 N1 N2 116.2285p
L3 N2 N3 57.7758p
L4 N3 N4 291.3934p
L5 N4 N5 76.1910p
L6 N5 N6 53.9027p
R1 2 N1 727.0696m
R2 2 N2 420.3238m
R3 2 N3 267.8926m
R4 2 N4 214.1069m
R5 2 N5 182.4512m
R6 2 N6 88.8345m
R7 2 N7 1.946
R8 2 1 1000000
.ends 0603_744761020A_2n
*******
.subckt 0603_744761033A_3.3n 1 2
C1 1 N7 0.228176204146948p
L1 1 N1 3.1n
L2 N1 N2 74.6789p
L3 N2 N3 54.4807p
L4 N3 N4 290.7303p
L5 N4 N5 76.1888p
L6 N5 N6 53.9010p
R1 2 N1 716.9716m
R2 2 N2 418.1686m
R3 2 N3 266.6832m
R4 2 N4 214.0411m
R5 2 N5 182.5034m
R6 2 N6 88.8381m
R7 2 N7 1.946
R8 2 1 1000000
.ends 0603_744761033A_3.3n
*******
.subckt 0603_744761036A_3.6n 1 2
C1 1 N7 0.202131386054143p
L1 1 N1 3.4n
L2 N1 N2 147.3304p
L3 N2 N3 36.2573p
L4 N3 N4 290.2187p
L5 N4 N5 76.2384p
L6 N5 N6 53.9414p
R1 2 N1 779.7842m
R2 2 N2 416.0625m
R3 2 N3 265.7198m
R4 2 N4 218.4858m
R5 2 N5 189.5536m
R6 2 N6 89.1102m
R7 2 N7 1.946
R8 2 1 1000000
.ends 0603_744761036A_3.6n
*******
.subckt 0603_744761039A_3.9n 1 2
C1 1 N7 0.180415219193454p
L1 1 N1 3.6n
L2 N1 N2 114.9991p
L3 N2 N3 172.8258p
L4 N3 N4 424.0175p
L5 N4 N5 77.1268p
L6 N5 N6 54.3887p
R1 2 N1 832.0440m
R2 2 N2 396.5298m
R3 2 N3 332.8480m
R4 2 N4 279.0579m
R5 2 N5 250.3686m
R6 2 N6 92.0094m
R7 2 N7 1.9461
R8 2 1 1000000
.ends 0603_744761039A_3.9n
*******
.subckt 0603_744761043A_4.3n 1 2
C1 1 N7 0.169226276696492p
L1 1 N1 4n
L2 N1 N2 122.8906p
L3 N2 N3 254.4246p
L4 N3 N4 522.8964p
L5 N4 N5 78.1133p
L6 N5 N6 55.0456p
R1 2 N1 1.3831
R2 2 N2 431.6943m
R3 2 N3 277.5790m
R4 2 N4 380.2072m
R5 2 N5 362.3595m
R6 2 N6 102.2510m
R7 2 N7 1.9462
R8 2 1 1000000
.ends 0603_744761043A_4.3n
*******
.subckt 0603_744761047A_4.7n 1 2
C1 1 N7 0.160208824188283p
L1 1 N1 4n
L2 N1 N2 133.4552p
L3 N2 N3 339.8837p
L4 N3 N4 550.3992p
L5 N4 N5 78.2267p
L6 N5 N6 55.0949p
R1 2 N1 1.3941
R2 2 N2 362.6733m
R3 2 N3 365.5944m
R4 2 N4 377.4310m
R5 2 N5 356.9140m
R6 2 N6 101.5009m
R7 2 N7 1.9462
R8 2 1 1000000
.ends 0603_744761047A_4.7n
*******
.subckt 0603_744761051A_5.1n 1 2
C1 1 N7 0.15286934003682p
L1 1 N1 4.5n
L2 N1 N2 135.5417p
L3 N2 N3 367.8063p
L4 N3 N4 569.0129p
L5 N4 N5 78.4327p
L6 N5 N6 55.2414p
R1 2 N1 1.3866
R2 2 N2 492.9421m
R3 2 N3 350.3851m
R4 2 N4 396.7967m
R5 2 N5 377.7113m
R6 2 N6 103.9987m
R7 2 N7 1.9462
R8 2 1 1000000
.ends 0603_744761051A_5.1n
*******
.subckt 0603_744761051GA_5.1n 1 2
C1 1 N7 0.15286934003682p
L1 1 N1 4.5n
L2 N1 N2 135.5417p
L3 N2 N3 367.8063p
L4 N3 N4 569.0129p
L5 N4 N5 78.4327p
L6 N5 N6 55.2414p
R1 2 N1 1.3866
R2 2 N2 492.9421m
R3 2 N3 350.3851m
R4 2 N4 396.7967m
R5 2 N5 377.7113m
R6 2 N6 103.9987m
R7 2 N7 1.9462
R8 2 1 1000000
.ends 0603_744761051GA_5.1n
*******
.subckt 0603_744761056A_5.6n 1 2
C1 1 N7 0.149529496899416p
L1 1 N1 4.85n
L2 N1 N2 199.3958p
L3 N2 N3 379.5339p
L4 N3 N4 699.3882p
L5 N4 N5 79.4612p
L6 N5 N6 55.9148p
R1 2 N1 1.5662
R2 2 N2 474.9501m
R3 2 N3 373.0310m
R4 2 N4 463.9700m
R5 2 N5 444.8165m
R6 2 N6 112.8385m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761056A_5.6n
*******
.subckt 0603_744761056GA_5.6n 1 2
C1 1 N7 0.149529496899416p
L1 1 N1 4.85n
L2 N1 N2 199.3958p
L3 N2 N3 379.5339p
L4 N3 N4 699.3882p
L5 N4 N5 79.4612p
L6 N5 N6 55.9148p
R1 2 N1 1.5662
R2 2 N2 474.9501m
R3 2 N3 373.0310m
R4 2 N4 463.9700m
R5 2 N5 444.8165m
R6 2 N6 112.8385m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761056GA_5.6n
*******
.subckt 0603_744761068A_6.8n 1 2
C1 1 N7 0.110732569659548p
L1 1 N1 6n
L2 N1 N2 147.5265p
L3 N2 N3 330.3889p
L4 N3 N4 703.1805p
L5 N4 N5 79.5071p
L6 N5 N6 55.9479p
R1 2 N1 1.5489
R2 2 N2 468.1799m
R3 2 N3 343.1308m
R4 2 N4 467.2763m
R5 2 N5 448.3296m
R6 2 N6 113.3581m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761068A_6.8n
*******
.subckt 0603_744761068GA_6.8n 1 2
C1 1 N7 0.110732569659548p
L1 1 N1 6n
L2 N1 N2 147.5265p
L3 N2 N3 330.3889p
L4 N3 N4 703.1805p
L5 N4 N5 79.5071p
L6 N5 N6 55.9479p
R1 2 N1 1.5489
R2 2 N2 468.1799m
R3 2 N3 343.1308m
R4 2 N4 467.2763m
R5 2 N5 448.3296m
R6 2 N6 113.3581m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761068GA_6.8n
*******
.subckt 0603_744761075A_7.5n 1 2
C1 1 N7 0.146587365594682p
L1 1 N1 7n
L2 N1 N2 266.3163p
L3 N2 N3 330.5894p
L4 N3 N4 703.0119p
L5 N4 N5 79.5084p
L6 N5 N6 55.9499p
R1 2 N1 1.559
R2 2 N2 480.3369m
R3 2 N3 340.9147m
R4 2 N4 467.4884m
R5 2 N5 448.5782m
R6 2 N6 113.3947m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761075A_7.5n
*******
.subckt 0603_744761075GA_7.5n 1 2
C1 1 N7 0.146587365594682p
L1 1 N1 7n
L2 N1 N2 266.3163p
L3 N2 N3 330.5894p
L4 N3 N4 703.0119p
L5 N4 N5 79.5084p
L6 N5 N6 55.9499p
R1 2 N1 1.559
R2 2 N2 480.3369m
R3 2 N3 340.9147m
R4 2 N4 467.4884m
R5 2 N5 448.5782m
R6 2 N6 113.3947m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761075GA_7.5n
*******
.subckt 0603_744761082A_8.2n 1 2
C1 1 N7 0.145985849824571p
L1 1 N1 7.5n
L2 N1 N2 204.8467p
L3 N2 N3 316.4480p
L4 N3 N4 694.5175p
L5 N4 N5 79.4764p
L6 N5 N6 55.9368p
R1 2 N1 1.6042
R2 2 N2 478.2306m
R3 2 N3 292.7134m
R4 2 N4 470.0855m
R5 2 N5 452.0271m
R6 2 N6 113.9566m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761082A_8.2n
*******
.subckt 0603_744761082GA_8.2n 1 2
C1 1 N7 0.145985849824571p
L1 1 N1 7.5n
L2 N1 N2 204.8467p
L3 N2 N3 316.4480p
L4 N3 N4 694.5175p
L5 N4 N5 79.4764p
L6 N5 N6 55.9368p
R1 2 N1 1.6042
R2 2 N2 478.2306m
R3 2 N3 292.7134m
R4 2 N4 470.0855m
R5 2 N5 452.0271m
R6 2 N6 113.9566m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761082GA_8.2n
*******
.subckt 0603_744761087A_8.7n 1 2
C1 1 N7 0.137595858455343p
L1 1 N1 8n
L2 N1 N2 183.9417p
L3 N2 N3 347.2170p
L4 N3 N4 698.0674p
L5 N4 N5 79.5063p
L6 N5 N6 55.9572p
R1 2 N1 1.5845
R2 2 N2 533.2879m
R3 2 N3 295.2036m
R4 2 N4 471.8835m
R5 2 N5 453.8292m
R6 2 N6 114.2213m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761087A_8.7n
*******
.subckt 0603_744761087GA_8.7n 1 2
C1 1 N7 0.137595858455343p
L1 1 N1 8n
L2 N1 N2 183.9417p
L3 N2 N3 347.2170p
L4 N3 N4 698.0674p
L5 N4 N5 79.5063p
L6 N5 N6 55.9572p
R1 2 N1 1.5845
R2 2 N2 533.2879m
R3 2 N3 295.2036m
R4 2 N4 471.8835m
R5 2 N5 453.8292m
R6 2 N6 114.2213m
R7 2 N7 1.9463
R8 2 1 1000000
.ends 0603_744761087GA_8.7n
*******
.subckt 0603_744761091A_9.1n 1 2
C1 1 N7 0.173971818507974p
L1 1 N1 8.3n
L2 N1 N2 205.5187p
L3 N2 N3 443.7610p
L4 N3 N4 782.5231p
L5 N4 N5 80.1794p
L6 N5 N6 56.4112p
R1 2 N1 1.86
R2 2 N2 563.5912m
R3 2 N3 346.8095m
R4 2 N4 512.6628m
R5 2 N5 494.2985m
R6 2 N6 120.3655m
R7 2 N7 1.9467
R8 2 1 1000000
.ends 0603_744761091A_9.1n
*******
.subckt 0603_744761091GA_9.1n 1 2
C1 1 N7 0.173971818507974p
L1 1 N1 8.3n
L2 N1 N2 205.5187p
L3 N2 N3 443.7610p
L4 N3 N4 782.5231p
L5 N4 N5 80.1794p
L6 N5 N6 56.4112p
R1 2 N1 1.86
R2 2 N2 563.5912m
R3 2 N3 346.8095m
R4 2 N4 512.6628m
R5 2 N5 494.2985m
R6 2 N6 120.3655m
R7 2 N7 1.9467
R8 2 1 1000000
.ends 0603_744761091GA_9.1n
*******
.subckt 0603_744761095A_9.5n 1 2
C1 1 N7 0.131671458218381p
L1 1 N1 8.7n
L2 N1 N2 253.7536p
L3 N2 N3 547.8332p
L4 N3 N4 760.5202p
L5 N4 N5 75.6049p
L6 N5 N6 53.7667p
R1 2 N1 2.4057
R2 2 N2 387.4905m
R3 2 N3 449.5366m
R4 2 N4 500.6298m
R5 2 N5 481.4257m
R6 2 N6 303.0031m
R7 2 N7 1.9468
R8 2 1 1000000
.ends 0603_744761095A_9.5n
*******
.subckt 0603_744761095GA_9.5n 1 2
C1 1 N7 0.131671458218381p
L1 1 N1 8.7n
L2 N1 N2 253.7536p
L3 N2 N3 547.8332p
L4 N3 N4 760.5202p
L5 N4 N5 75.6049p
L6 N5 N6 53.7667p
R1 2 N1 2.4057
R2 2 N2 387.4905m
R3 2 N3 449.5366m
R4 2 N4 500.6298m
R5 2 N5 481.4257m
R6 2 N6 303.0031m
R7 2 N7 1.9468
R8 2 1 1000000
.ends 0603_744761095GA_9.5n
*******
.subckt 0603_744761110A_10n 1 2
C1 1 N7 0.109940524196011p
L1 1 N1 9.5n
L2 N1 N2 258.8631p
L3 N2 N3 608.4738p
L4 N3 N4 775.7247p
L5 N4 N5 75.6980p
L6 N5 N6 53.8050p
R1 2 N1 2.4586
R2 2 N2 625.4426m
R3 2 N3 468.3310m
R4 2 N4 515.5851m
R5 2 N5 496.6291m
R6 2 N6 338.5348m
R7 2 N7 1.9469
R8 2 1 1000000
.ends 0603_744761110A_10n
*******
.subckt 0603_744761110GA_10n 1 2
C1 1 N7 0.109940524196011p
L1 1 N1 9.5n
L2 N1 N2 258.8631p
L3 N2 N3 608.4738p
L4 N3 N4 775.7247p
L5 N4 N5 75.6980p
L6 N5 N6 53.8050p
R1 2 N1 2.4586
R2 2 N2 625.4426m
R3 2 N3 468.3310m
R4 2 N4 515.5851m
R5 2 N5 496.6291m
R6 2 N6 338.5348m
R7 2 N7 1.9469
R8 2 1 1000000
.ends 0603_744761110GA_10n
*******
.subckt 0603_744761111A_11n 1 2
C1 1 N7 0.143922140765687p
L1 1 N1 10.5n
L2 N1 N2 155.4961p
L3 N2 N3 444.5546p
L4 N3 N4 750.7819p
L5 N4 N5 75.1470p
L6 N5 N6 53.5356p
R1 2 N1 2.4439
R2 2 N2 756.4287m
R3 2 N3 301.4124m
R4 2 N4 507.2606m
R5 2 N5 490.0777m
R6 2 N6 330.2335m
R7 2 N7 1.937
R8 2 1 1000000
.ends 0603_744761111A_11n
*******
.subckt 0603_744761111GA_11n 1 2
C1 1 N7 0.143922140765687p
L1 1 N1 10.5n
L2 N1 N2 155.4961p
L3 N2 N3 444.5546p
L4 N3 N4 750.7819p
L5 N4 N5 75.1470p
L6 N5 N6 53.5356p
R1 2 N1 2.4439
R2 2 N2 756.4287m
R3 2 N3 301.4124m
R4 2 N4 507.2606m
R5 2 N5 490.0777m
R6 2 N6 330.2335m
R7 2 N7 1.937
R8 2 1 1000000
.ends 0603_744761111GA_11n
*******
.subckt 0603_744761112A_12n 1 2
C1 1 N7 0.131928629035214p
L1 1 N1 11.5n
L2 N1 N2 233.6059p
L3 N2 N3 508.6165p
L4 N3 N4 831.9102p
L5 N4 N5 75.6267p
L6 N5 N6 53.7413p
R1 2 N1 2.4187
R2 2 N2 928.7942m
R3 2 N3 433.9025m
R4 2 N4 552.9997m
R5 2 N5 534.0380m
R6 2 N6 413.0624m
R7 2 N7 1.9294
R8 2 1 1000000
.ends 0603_744761112A_12n
*******
.subckt 0603_744761112GA_12n 1 2
C1 1 N7 0.131928629035214p
L1 1 N1 11.5n
L2 N1 N2 233.6059p
L3 N2 N3 508.6165p
L4 N3 N4 831.9102p
L5 N4 N5 75.6267p
L6 N5 N6 53.7413p
R1 2 N1 2.4187
R2 2 N2 928.7942m
R3 2 N3 433.9025m
R4 2 N4 552.9997m
R5 2 N5 534.0380m
R6 2 N6 413.0624m
R7 2 N7 1.9294
R8 2 1 1000000
.ends 0603_744761112GA_12n
*******
.subckt 0603_744761113A_13n 1 2
C1 1 N7 0.121780272955582p
L1 1 N1 12.5n
L2 N1 N2 201.8003p
L3 N2 N3 502.9679p
L4 N3 N4 831.9408p
L5 N4 N5 75.6264p
L6 N5 N6 53.7402p
R1 2 N1 2.4176
R2 2 N2 922.1835m
R3 2 N3 432.0556m
R4 2 N4 553.0946m
R5 2 N5 534.1373m
R6 2 N6 413.2267m
R7 2 N7 1.9293
R8 2 1 1000000
.ends 0603_744761113A_13n
*******
.subckt 0603_744761113GA_13n 1 2
C1 1 N7 0.121780272955582p
L1 1 N1 12.5n
L2 N1 N2 201.8003p
L3 N2 N3 502.9679p
L4 N3 N4 831.9408p
L5 N4 N5 75.6264p
L6 N5 N6 53.7402p
R1 2 N1 2.4176
R2 2 N2 922.1835m
R3 2 N3 432.0556m
R4 2 N4 553.0946m
R5 2 N5 534.1373m
R6 2 N6 413.2267m
R7 2 N7 1.9293
R8 2 1 1000000
.ends 0603_744761113GA_13n
*******
.subckt 0603_744761115A_15n 1 2
C1 1 N7 0.105542903228171p
L1 1 N1 14.3n
L2 N1 N2 338.6149p
L3 N2 N3 619.0164p
L4 N3 N4 934.6943p
L5 N4 N5 76.1373p
L6 N5 N6 53.9019p
R1 2 N1 2.435
R2 2 N2 925.4044m
R3 2 N3 603.5517m
R4 2 N4 600.2547m
R5 2 N5 578.6399m
R6 2 N6 479.7717m
R7 2 N7 1.9331
R8 2 1 1000000
.ends 0603_744761115A_15n
*******
.subckt 0603_744761115GA_15n 1 2
C1 1 N7 0.105542903228171p
L1 1 N1 14.3n
L2 N1 N2 338.6149p
L3 N2 N3 619.0164p
L4 N3 N4 934.6943p
L5 N4 N5 76.1373p
L6 N5 N6 53.9019p
R1 2 N1 2.435
R2 2 N2 925.4044m
R3 2 N3 603.5517m
R4 2 N4 600.2547m
R5 2 N5 578.6399m
R6 2 N6 479.7717m
R7 2 N7 1.9331
R8 2 1 1000000
.ends 0603_744761115GA_15n
*******
.subckt 0603_744761116A_16n 1 2
C1 1 N7 0.145375899763321p
L1 1 N1 15.2n
L2 N1 N2 375.4590p
L3 N2 N3 710.9366p
L4 N3 N4 1.0513n
L5 N4 N5 76.7287p
L6 N5 N6 54.0824p
R1 2 N1 2.3999
R2 2 N2 1.031
R3 2 N3 707.3204m
R4 2 N4 669.5653m
R5 2 N5 646.5994m
R6 2 N6 570.8999m
R7 2 N7 1.9226
R8 2 1 1000000
.ends 0603_744761116A_16n
*******
.subckt 0603_744761116GA_16n 1 2
C1 1 N7 0.145375899763321p
L1 1 N1 15.2n
L2 N1 N2 375.4590p
L3 N2 N3 710.9366p
L4 N3 N4 1.0513n
L5 N4 N5 76.7287p
L6 N5 N6 54.0824p
R1 2 N1 2.3999
R2 2 N2 1.031
R3 2 N3 707.3204m
R4 2 N4 669.5653m
R5 2 N5 646.5994m
R6 2 N6 570.8999m
R7 2 N7 1.9226
R8 2 1 1000000
.ends 0603_744761116GA_16n
*******
.subckt 0603_744761118A_18n 1 2
C1 1 N7 0.146434829314146p
L1 1 N1 17.2n
L2 N1 N2 252.3963p
L3 N2 N3 738.6997p
L4 N3 N4 1.1678n
L5 N4 N5 77.3518p
L6 N5 N6 54.2682p
R1 2 N1 2.2938
R2 2 N2 1.4697
R3 2 N3 728.5670m
R4 2 N4 774.4066m
R5 2 N5 752.7530m
R6 2 N6 699.7297m
R7 2 N7 1.8424
R8 2 1 1000000
.ends 0603_744761118A_18n
*******
.subckt 0603_744761118GA_18n 1 2
C1 1 N7 0.146434829314146p
L1 1 N1 17.2n
L2 N1 N2 252.3963p
L3 N2 N3 738.6997p
L4 N3 N4 1.1678n
L5 N4 N5 77.3518p
L6 N5 N6 54.2682p
R1 2 N1 2.2938
R2 2 N2 1.4697
R3 2 N3 728.5670m
R4 2 N4 774.4066m
R5 2 N5 752.7530m
R6 2 N6 699.7297m
R7 2 N7 1.8424
R8 2 1 1000000
.ends 0603_744761118GA_18n
*******
.subckt 0603_744761120A_20n 1 2
C1 1 N7 0.140723870970894p
L1 1 N1 19n
L2 N1 N2 312.6360p
L3 N2 N3 738.4750p
L4 N3 N4 1.1676n
L5 N4 N5 77.3527p
L6 N5 N6 54.2699p
R1 2 N1 2.3006
R2 2 N2 1.4782
R3 2 N3 726.7858m
R4 2 N4 774.4871m
R5 2 N5 752.8442m
R6 2 N6 699.8346m
R7 2 N7 1.8431
R8 2 1 1000000
.ends 0603_744761120A_20n
*******
.subckt 0603_744761120GA_20n 1 2
C1 1 N7 0.140723870970894p
L1 1 N1 19n
L2 N1 N2 312.6360p
L3 N2 N3 738.4750p
L4 N3 N4 1.1676n
L5 N4 N5 77.3527p
L6 N5 N6 54.2699p
R1 2 N1 2.3006
R2 2 N2 1.4782
R3 2 N3 726.7858m
R4 2 N4 774.4871m
R5 2 N5 752.8442m
R6 2 N6 699.8346m
R7 2 N7 1.8431
R8 2 1 1000000
.ends 0603_744761120GA_20n
*******
.subckt 0603_744761122A_22n 1 2
C1 1 N7 0.127930791791722p
L1 1 N1 21n
L2 N1 N2 523.9604p
L3 N2 N3 701.2403p
L4 N3 N4 1.2497n
L5 N4 N5 77.7499p
L6 N5 N6 54.3800p
R1 2 N1 2.5051
R2 2 N2 1.4063
R3 2 N3 814.1749m
R4 2 N4 821.0948m
R5 2 N5 798.4407m
R6 2 N6 750.5338m
R7 2 N7 1.889
R8 2 1 1000000
.ends 0603_744761122A_22n
*******
.subckt 0603_744761122GA_22n 1 2
C1 1 N7 0.127930791791722p
L1 1 N1 21n
L2 N1 N2 523.9604p
L3 N2 N3 701.2403p
L4 N3 N4 1.2497n
L5 N4 N5 77.7499p
L6 N5 N6 54.3800p
R1 2 N1 2.5051
R2 2 N2 1.4063
R3 2 N3 814.1749m
R4 2 N4 821.0948m
R5 2 N5 798.4407m
R6 2 N6 750.5338m
R7 2 N7 1.889
R8 2 1 1000000
.ends 0603_744761122GA_22n
*******
.subckt 0603_744761124A_24n 1 2
C1 1 N7 0.156128555071259p
L1 1 N1 23n
L2 N1 N2 422.6565p
L3 N2 N3 856.9138p
L4 N3 N4 1.4168n
L5 N4 N5 78.5752p
L6 N5 N6 54.6163p
R1 2 N1 2.2819
R2 2 N2 1.5684
R3 2 N3 939.0760m
R4 2 N4 909.0252m
R5 2 N5 884.2852m
R6 2 N6 843.7675m
R7 2 N7 1.7593
R8 2 1 1000000
.ends 0603_744761124A_24n
*******
.subckt 0603_744761124GA_24n 1 2
C1 1 N7 0.156128555071259p
L1 1 N1 23n
L2 N1 N2 422.6565p
L3 N2 N3 856.9138p
L4 N3 N4 1.4168n
L5 N4 N5 78.5752p
L6 N5 N6 54.6163p
R1 2 N1 2.2819
R2 2 N2 1.5684
R3 2 N3 939.0760m
R4 2 N4 909.0252m
R5 2 N5 884.2852m
R6 2 N6 843.7675m
R7 2 N7 1.7593
R8 2 1 1000000
.ends 0603_744761124GA_24n
*******
.subckt 0603_744761127A_27n 1 2
C1 1 N7 0.119663155587495p
L1 1 N1 25.5n
L2 N1 N2 551.5124p
L3 N2 N3 615.4934p
L4 N3 N4 1.4153n
L5 N4 N5 78.5859p
L6 N5 N6 54.6175p
R1 2 N1 2.5631
R2 2 N2 1.398
R3 2 N3 862.0667m
R4 2 N4 915.6808m
R5 2 N5 891.3432m
R6 2 N6 851.4592m
R7 2 N7 1.8232
R8 2 1 1000000
.ends 0603_744761127A_27n
*******
.subckt 0603_744761127GA_27n 1 2
C1 1 N7 0.119663155587495p
L1 1 N1 25.5n
L2 N1 N2 551.5124p
L3 N2 N3 615.4934p
L4 N3 N4 1.4153n
L5 N4 N5 78.5859p
L6 N5 N6 54.6175p
R1 2 N1 2.5631
R2 2 N2 1.398
R3 2 N3 862.0667m
R4 2 N4 915.6808m
R5 2 N5 891.3432m
R6 2 N6 851.4592m
R7 2 N7 1.8232
R8 2 1 1000000
.ends 0603_744761127GA_27n
*******
.subckt 0603_744761130A_30n 1 2
C1 1 N7 0.135094916132059p
L1 1 N1 28.5n
L2 N1 N2 712.0090p
L3 N2 N3 980.9304p
L4 N3 N4 1.7527n
L5 N4 N5 80.1498p
L6 N5 N6 55.0280p
R1 2 N1 3.1033
R2 2 N2 1.2438
R3 2 N3 1.3515
R4 2 N4 1.0781
R5 2 N5 1.0499
R6 2 N6 1.0187
R7 2 N7 2.0312
R8 2 1 1000000
.ends 0603_744761130A_30n
*******
.subckt 0603_744761130GA_30n 1 2
C1 1 N7 0.135094916132059p
L1 1 N1 28.5n
L2 N1 N2 712.0090p
L3 N2 N3 980.9304p
L4 N3 N4 1.7527n
L5 N4 N5 80.1498p
L6 N5 N6 55.0280p
R1 2 N1 3.1033
R2 2 N2 1.2438
R3 2 N3 1.3515
R4 2 N4 1.0781
R5 2 N5 1.0499
R6 2 N6 1.0187
R7 2 N7 2.0312
R8 2 1 1000000
.ends 0603_744761130GA_30n
*******
.subckt 0603_744761133A_33n 1 2
C1 1 N7 0.145101087098362p
L1 1 N1 31.5n
L2 N1 N2 628.7195p
L3 N2 N3 758.2566p
L4 N3 N4 1.9073n
L5 N4 N5 82.9611p
L6 N5 N6 58.0554p
R1 2 N1 2.226
R2 2 N2 1.8845
R3 2 N3 784.2121m
R4 2 N4 1.0094
R5 2 N5 970.9148m
R6 2 N6 930.9504m
R7 2 N7 3.6753
R8 2 1 1000000
.ends 0603_744761133A_33n
*******
.subckt 0603_744761133GA_33n 1 2
C1 1 N7 0.145101087098362p
L1 1 N1 31.5n
L2 N1 N2 628.7195p
L3 N2 N3 758.2566p
L4 N3 N4 1.9073n
L5 N4 N5 82.9611p
L6 N5 N6 58.0554p
R1 2 N1 2.226
R2 2 N2 1.8845
R3 2 N3 784.2121m
R4 2 N4 1.0094
R5 2 N5 970.9148m
R6 2 N6 930.9504m
R7 2 N7 3.6753
R8 2 1 1000000
.ends 0603_744761133GA_33n
*******
.subckt 0603_744761136A_36n 1 2
C1 1 N7 0.133009329840165p
L1 1 N1 34n
L2 N1 N2 845.8858p
L3 N2 N3 618.5224p
L4 N3 N4 2.2849n
L5 N4 N5 87.3132p
L6 N5 N6 62.1356p
R1 2 N1 2.8675
R2 2 N2 1.9258
R3 2 N3 1.1584
R4 2 N4 1.122
R5 2 N5 1.0779
R6 2 N6 1.0404
R7 2 N7 4.7014
R8 2 1 1000000
.ends 0603_744761136A_36n
*******
.subckt 0603_744761136GA_36n 1 2
C1 1 N7 0.133009329840165p
L1 1 N1 34n
L2 N1 N2 845.8858p
L3 N2 N3 618.5224p
L4 N3 N4 2.2849n
L5 N4 N5 87.3132p
L6 N5 N6 62.1356p
R1 2 N1 2.8675
R2 2 N2 1.9258
R3 2 N3 1.1584
R4 2 N4 1.122
R5 2 N5 1.0779
R6 2 N6 1.0404
R7 2 N7 4.7014
R8 2 1 1000000
.ends 0603_744761136GA_36n
*******
.subckt 0603_744761139A_39n 1 2
C1 1 N7 0.134193138243065p
L1 1 N1 37n
L2 N1 N2 1.0775n
L3 N2 N3 654.9051p
L4 N3 N4 3.2695n
L5 N4 N5 75.6328p
L6 N5 N6 54.0106p
R1 2 N1 2.6838
R2 2 N2 2.0236
R3 2 N3 1.3041
R4 2 N4 1.3015
R5 2 N5 1.2694
R6 2 N6 1.2431
R7 2 N7 6.188
R8 2 1 1000000
.ends 0603_744761139A_39n
*******
.subckt 0603_744761139GA_39n 1 2
C1 1 N7 0.134193138243065p
L1 1 N1 37n
L2 N1 N2 1.0775n
L3 N2 N3 654.9051p
L4 N3 N4 3.2695n
L5 N4 N5 75.6328p
L6 N5 N6 54.0106p
R1 2 N1 2.6838
R2 2 N2 2.0236
R3 2 N3 1.3041
R4 2 N4 1.3015
R5 2 N5 1.2694
R6 2 N6 1.2431
R7 2 N7 6.188
R8 2 1 1000000
.ends 0603_744761139GA_39n
*******
.subckt 0603_744761143A_43n 1 2
C1 1 N7 0.147269167295122p
L1 1 N1 40.7n
L2 N1 N2 1.5208n
L3 N2 N3 429.8598p
L4 N3 N4 5.5588n
L5 N4 N5 83.8588p
L6 N5 N6 65.3852p
R1 2 N1 2.3283
R2 2 N2 2.1462
R3 2 N3 1.4653
R4 2 N4 1.5709
R5 2 N5 1.5485
R6 2 N6 1.5306
R7 2 N7 7.5346
R8 2 1 1000000
.ends 0603_744761143A_43n
*******
.subckt 0603_744761143GA_43n 1 2
C1 1 N7 0.147269167295122p
L1 1 N1 40.7n
L2 N1 N2 1.5208n
L3 N2 N3 429.8598p
L4 N3 N4 5.5588n
L5 N4 N5 83.8588p
L6 N5 N6 65.3852p
R1 2 N1 2.3283
R2 2 N2 2.1462
R3 2 N3 1.4653
R4 2 N4 1.5709
R5 2 N5 1.5485
R6 2 N6 1.5306
R7 2 N7 7.5346
R8 2 1 1000000
.ends 0603_744761143GA_43n
*******
.subckt 0603_744761147A_47n 1 2
C1 1 N7 0.134735621142346p
L1 1 N1 44.5n
L2 N1 N2 1.3981n
L3 N2 N3 681.0799p
L4 N3 N4 3.1208n
L5 N4 N5 90.6030p
L6 N5 N6 74.0832p
R1 2 N1 3.2669
R2 2 N2 2.2164
R3 2 N3 1.5398
R4 2 N4 1.2718
R5 2 N5 1.2385
R6 2 N6 1.2113
R7 2 N7 9.9034
R8 2 1 1000000
.ends 0603_744761147A_47n
*******
.subckt 0603_744761147GA_47n 1 2
C1 1 N7 0.134735621142346p
L1 1 N1 44.5n
L2 N1 N2 1.3981n
L3 N2 N3 681.0799p
L4 N3 N4 3.1208n
L5 N4 N5 90.6030p
L6 N5 N6 74.0832p
R1 2 N1 3.2669
R2 2 N2 2.2164
R3 2 N3 1.5398
R4 2 N4 1.2718
R5 2 N5 1.2385
R6 2 N6 1.2113
R7 2 N7 9.9034
R8 2 1 1000000
.ends 0603_744761147GA_47n
*******
.subckt 0603_744761151A_51n 1 2
C1 1 N7 0.137582406033138p
L1 1 N1 49n
L2 N1 N2 1.7938n
L3 N2 N3 61.2233p
L4 N3 N4 4.8127n
L5 N4 N5 91.0957p
L6 N5 N6 74.4174p
R1 2 N1 3.7335
R2 2 N2 2.3161
R3 2 N3 1.5603
R4 2 N4 1.1437
R5 2 N5 1.1004
R6 2 N6 1.0651
R7 2 N7 7.8229
R8 2 1 1000000
.ends 0603_744761151A_51n
*******
.subckt 0603_744761151GA_51n 1 2
C1 1 N7 0.137582406033138p
L1 1 N1 49n
L2 N1 N2 1.7938n
L3 N2 N3 61.2233p
L4 N3 N4 4.8127n
L5 N4 N5 91.0957p
L6 N5 N6 74.4174p
R1 2 N1 3.7335
R2 2 N2 2.3161
R3 2 N3 1.5603
R4 2 N4 1.1437
R5 2 N5 1.1004
R6 2 N6 1.0651
R7 2 N7 7.8229
R8 2 1 1000000
.ends 0603_744761151GA_51n
*******
.subckt 0603_744761156A_56n 1 2
C1 1 N7 0.125298262637322p
L1 1 N1 53.5n
L2 N1 N2 2.0122n
L3 N2 N3 275.1924p
L4 N3 N4 5.3841n
L5 N4 N5 91.8945p
L6 N5 N6 75.3308p
R1 2 N1 3.2927
R2 2 N2 2.432
R3 2 N3 1.7796
R4 2 N4 1.4663
R5 2 N5 1.4413
R6 2 N6 1.4221
R7 2 N7 6.4387
R8 2 1 1000000
.ends 0603_744761156A_56n
*******
.subckt 0603_744761156GA_56n 1 2
C1 1 N7 0.125298262637322p
L1 1 N1 53.5n
L2 N1 N2 2.0122n
L3 N2 N3 275.1924p
L4 N3 N4 5.3841n
L5 N4 N5 91.8945p
L6 N5 N6 75.3308p
R1 2 N1 3.2927
R2 2 N2 2.432
R3 2 N3 1.7796
R4 2 N4 1.4663
R5 2 N5 1.4413
R6 2 N6 1.4221
R7 2 N7 6.4387
R8 2 1 1000000
.ends 0603_744761156GA_56n
*******
.subckt 0603_744761162A_62n 1 2
C1 1 N7 0.14136788020293p
L1 1 N1 59n
L2 N1 N2 1.8430n
L3 N2 N3 1.1817n
L4 N3 N4 4.8336n
L5 N4 N5 75.3806p
L6 N5 N6 53.6520p
R1 2 N1 4.1464
R2 2 N2 2.1423
R3 2 N3 1.606
R4 2 N4 1.1632
R5 2 N5 1.1216
R6 2 N6 1.0869
R7 2 N7 5.1102
R8 2 1 1000000
.ends 0603_744761162A_62n
*******
.subckt 0603_744761162GA_62n 1 2
C1 1 N7 0.14136788020293p
L1 1 N1 59n
L2 N1 N2 1.8430n
L3 N2 N3 1.1817n
L4 N3 N4 4.8336n
L5 N4 N5 75.3806p
L6 N5 N6 53.6520p
R1 2 N1 4.1464
R2 2 N2 2.1423
R3 2 N3 1.606
R4 2 N4 1.1632
R5 2 N5 1.1216
R6 2 N6 1.0869
R7 2 N7 5.1102
R8 2 1 1000000
.ends 0603_744761162GA_62n
*******
.subckt 0603_744761168A_68n 1 2
C1 1 N7 0.128894243714436p
L1 1 N1 65n
L2 N1 N2 1.9806n
L3 N2 N3 1.4057n
L4 N3 N4 5.2311n
L5 N4 N5 75.7141p
L6 N5 N6 54.0801p
R1 2 N1 4.6712
R2 2 N2 2.3348
R3 2 N3 1.9478
R4 2 N4 1.3003
R5 2 N5 1.2676
R6 2 N6 1.2411
R7 2 N7 5.2558
R8 2 1 1000000
.ends 0603_744761168A_68n
*******
.subckt 0603_744761168GA_68n 1 2
C1 1 N7 0.128894243714436p
L1 1 N1 65n
L2 N1 N2 1.9806n
L3 N2 N3 1.4057n
L4 N3 N4 5.2311n
L5 N4 N5 75.7141p
L6 N5 N6 54.0801p
R1 2 N1 4.6712
R2 2 N2 2.3348
R3 2 N3 1.9478
R4 2 N4 1.3003
R5 2 N5 1.2676
R6 2 N6 1.2411
R7 2 N7 5.2558
R8 2 1 1000000
.ends 0603_744761168GA_68n
*******
.subckt 0603_744761172A_72n 1 2
C1 1 N7 0.121733452396967p
L1 1 N1 68n
L2 N1 N2 2.3382n
L3 N2 N3 1.4425n
L4 N3 N4 6.9996n
L5 N4 N5 79.7514p
L6 N5 N6 59.5651p
R1 2 N1 4.3456
R2 2 N2 2.6681
R3 2 N3 2.6651
R4 2 N4 2.2368
R5 2 N5 2.2355
R6 2 N6 2.2352
R7 2 N7 4.0353
R8 2 1 1000000
.ends 0603_744761172A_72n
*******
.subckt 0603_744761172GA_72n 1 2
C1 1 N7 0.121733452396967p
L1 1 N1 68n
L2 N1 N2 2.3382n
L3 N2 N3 1.4425n
L4 N3 N4 6.9996n
L5 N4 N5 79.7514p
L6 N5 N6 59.5651p
R1 2 N1 4.3456
R2 2 N2 2.6681
R3 2 N3 2.6651
R4 2 N4 2.2368
R5 2 N5 2.2355
R6 2 N6 2.2352
R7 2 N7 4.0353
R8 2 1 1000000
.ends 0603_744761172GA_72n
*******
.subckt 0603_744761182A_82n 1 2
C1 1 N7 0.106887909421728p
L1 1 N1 78n
L2 N1 N2 1.9181n
L3 N2 N3 1.8685n
L4 N3 N4 4.6703n
L5 N4 N5 78.3642p
L6 N5 N6 57.7653p
R1 2 N1 9.1611
R2 2 N2 3.1169
R3 2 N3 3.5069
R4 2 N4 2.3056
R5 2 N5 2.3045
R6 2 N6 2.3043
R7 2 N7 6.5091
R8 2 1 1000000
.ends 0603_744761182A_82n
*******
.subckt 0603_744761182GA_82n 1 2
C1 1 N7 0.106887909421728p
L1 1 N1 78n
L2 N1 N2 1.9181n
L3 N2 N3 1.8685n
L4 N3 N4 4.6703n
L5 N4 N5 78.3642p
L6 N5 N6 57.7653p
R1 2 N1 9.1611
R2 2 N2 3.1169
R3 2 N3 3.5069
R4 2 N4 2.3056
R5 2 N5 2.3045
R6 2 N6 2.3043
R7 2 N7 6.5091
R8 2 1 1000000
.ends 0603_744761182GA_82n
*******
.subckt 0603_744761190A_90n 1 2
C1 1 N7 0.097386761917574p
L1 1 N1 85n
L2 N1 N2 2.1649n
L3 N2 N3 1.9138n
L4 N3 N4 5.4017n
L5 N4 N5 78.3693p
L6 N5 N6 57.7377p
R1 2 N1 9.1716
R2 2 N2 3.1994
R3 2 N3 3.5239
R4 2 N4 2.3071
R5 2 N5 2.3059
R6 2 N6 2.3056
R7 2 N7 6.5051
R8 2 1 1000000
.ends 0603_744761190A_90n
*******
.subckt 0603_744761190GA_90n 1 2
C1 1 N7 0.097386761917574p
L1 1 N1 85n
L2 N1 N2 2.1649n
L3 N2 N3 1.9138n
L4 N3 N4 5.4017n
L5 N4 N5 78.3693p
L6 N5 N6 57.7377p
R1 2 N1 9.1716
R2 2 N2 3.1994
R3 2 N3 3.5239
R4 2 N4 2.3071
R5 2 N5 2.3059
R6 2 N6 2.3056
R7 2 N7 6.5051
R8 2 1 1000000
.ends 0603_744761190GA_90n
*******
.subckt 0603_744761210A_100n 1 2
C1 1 N7 0.129236208034495p
L1 1 N1 95n
L2 N1 N2 1.7596n
L3 N2 N3 2.6599n
L4 N3 N4 4.8152n
L5 N4 N5 79.7290p
L6 N5 N6 59.4010p
R1 2 N1 8.6434
R2 2 N2 4.4934
R3 2 N3 3.0072
R4 2 N4 2.4307
R5 2 N5 2.4294
R6 2 N6 2.429
R7 2 N7 8.7665
R8 2 1 1000000
.ends 0603_744761210A_100n
*******
.subckt 0603_744761210GA_100n 1 2
C1 1 N7 0.129236208034495p
L1 1 N1 95n
L2 N1 N2 1.7596n
L3 N2 N3 2.6599n
L4 N3 N4 4.8152n
L5 N4 N5 79.7290p
L6 N5 N6 59.4010p
R1 2 N1 8.6434
R2 2 N2 4.4934
R3 2 N3 3.0072
R4 2 N4 2.4307
R5 2 N5 2.4294
R6 2 N6 2.429
R7 2 N7 8.7665
R8 2 1 1000000
.ends 0603_744761210GA_100n
*******
.subckt 0603_744761211A_110n 1 2
C1 1 N7 0.117487461849541p
L1 1 N1 103n
L2 N1 N2 2.5532n
L3 N2 N3 2.6723n
L4 N3 N4 7.9368n
L5 N4 N5 81.0717p
L6 N5 N6 60.7542p
R1 2 N1 9.812
R2 2 N2 4.7682
R3 2 N3 2.544
R4 2 N4 3.1218
R5 2 N5 3.1203
R6 2 N6 3.1197
R7 2 N7 15.8764
R8 2 1 1000000
.ends 0603_744761211A_110n
*******
.subckt 0603_744761211GA_110n 1 2
C1 1 N7 0.117487461849541p
L1 1 N1 103n
L2 N1 N2 2.5532n
L3 N2 N3 2.6723n
L4 N3 N4 7.9368n
L5 N4 N5 81.0717p
L6 N5 N6 60.7542p
R1 2 N1 9.812
R2 2 N2 4.7682
R3 2 N3 2.544
R4 2 N4 3.1218
R5 2 N5 3.1203
R6 2 N6 3.1197
R7 2 N7 15.8764
R8 2 1 1000000
.ends 0603_744761211GA_110n
*******
.subckt 0603_744761212A_120n 1 2
C1 1 N7 0.124902844057007p
L1 1 N1 110n
L2 N1 N2 1.7582n
L3 N2 N3 4.6277n
L4 N3 N4 6.2084n
L5 N4 N5 81.0874p
L6 N5 N6 60.8523p
R1 2 N1 9.7768
R2 2 N2 5.0911
R3 2 N3 2.3746
R4 2 N4 3.1324
R5 2 N5 3.1311
R6 2 N6 3.1305
R7 2 N7 15.4321
R8 2 1 1000000
.ends 0603_744761212A_120n
*******
.subckt 0603_744761212GA_120n 1 2
C1 1 N7 0.124902844057007p
L1 1 N1 110n
L2 N1 N2 1.7582n
L3 N2 N3 4.6277n
L4 N3 N4 6.2084n
L5 N4 N5 81.0874p
L6 N5 N6 60.8523p
R1 2 N1 9.7768
R2 2 N2 5.0911
R3 2 N3 2.3746
R4 2 N4 3.1324
R5 2 N5 3.1311
R6 2 N6 3.1305
R7 2 N7 15.4321
R8 2 1 1000000
.ends 0603_744761212GA_120n
*******
.subckt 0603_744761215A_150n 1 2
C1 1 N7 75.2921f
L1 1 N1 140n
L2 N1 N2 4.8362n
L3 N2 N3 3.7158n
L4 N3 N4 13.6515n
L5 N4 N5 96.9943p
L6 N5 N6 81.7564p
R1 2 N1 9.7086
R2 2 N2 6.1901
R3 2 N3 2.4115
R4 2 N4 3.3958
R5 2 N5 3.3941
R6 2 N6 3.3934
R7 2 N7 36.0558
R8 2 1 1000000
.ends 0603_744761215A_150n
*******
.subckt 0603_744761215GA_150n 1 2
C1 1 N7 75.2921f
L1 1 N1 140n
L2 N1 N2 4.8362n
L3 N2 N3 3.7158n
L4 N3 N4 13.6515n
L5 N4 N5 96.9943p
L6 N5 N6 81.7564p
R1 2 N1 9.7086
R2 2 N2 6.1901
R3 2 N3 2.4115
R4 2 N4 3.3958
R5 2 N5 3.3941
R6 2 N6 3.3934
R7 2 N7 36.0558
R8 2 1 1000000
.ends 0603_744761215GA_150n
*******
.subckt 0603_744761216A_160n 1 2
C1 1 N7 85.3481f
L1 1 N1 150n
L2 N1 N2 4.7796n
L3 N2 N3 3.7524n
L4 N3 N4 14.0693n
L5 N4 N5 97.0075p
L6 N5 N6 81.7539p
R1 2 N1 9.7527
R2 2 N2 6.1887
R3 2 N3 2.4724
R4 2 N4 3.4069
R5 2 N5 3.4051
R6 2 N6 3.4044
R7 2 N7 38.8692
R8 2 1 1000000
.ends 0603_744761216A_160n
*******
.subckt 0603_744761216GA_160n 1 2
C1 1 N7 85.3481f
L1 1 N1 150n
L2 N1 N2 4.7796n
L3 N2 N3 3.7524n
L4 N3 N4 14.0693n
L5 N4 N5 97.0075p
L6 N5 N6 81.7539p
R1 2 N1 9.7527
R2 2 N2 6.1887
R3 2 N3 2.4724
R4 2 N4 3.4069
R5 2 N5 3.4051
R6 2 N6 3.4044
R7 2 N7 38.8692
R8 2 1 1000000
.ends 0603_744761216GA_160n
*******
.subckt 0603_744761218A_180n 1 2
C1 1 N7 85.7069f
L1 1 N1 168n
L2 N1 N2 5.8838n
L3 N2 N3 4.2359n
L4 N3 N4 15.1133n
L5 N4 N5 97.2459p
L6 N5 N6 81.9931p
R1 2 N1 9.8151
R2 2 N2 6.1909
R3 2 N3 2.5702
R4 2 N4 3.4249
R5 2 N5 3.423
R6 2 N6 3.4222
R7 2 N7 41.5186
R8 2 1 1000000
.ends 0603_744761218A_180n
*******
.subckt 0603_744761218GA_180n 1 2
C1 1 N7 85.7069f
L1 1 N1 168n
L2 N1 N2 5.8838n
L3 N2 N3 4.2359n
L4 N3 N4 15.1133n
L5 N4 N5 97.2459p
L6 N5 N6 81.9931p
R1 2 N1 9.8151
R2 2 N2 6.1909
R3 2 N3 2.5702
R4 2 N4 3.4249
R5 2 N5 3.423
R6 2 N6 3.4222
R7 2 N7 41.5186
R8 2 1 1000000
.ends 0603_744761218GA_180n
*******
.subckt 0603_744761220A_200n 1 2
C1 1 N7 96.5504f
L1 1 N1 185n
L2 N1 N2 7.0859n
L3 N2 N3 4.0485n
L4 N3 N4 19.1761n
L5 N4 N5 97.5419p
L6 N5 N6 82.1736p
R1 2 N1 9.9312
R2 2 N2 6.1986
R3 2 N3 2.8562
R4 2 N4 3.5033
R5 2 N5 3.501
R6 2 N6 3.5
R7 2 N7 41.8699
R8 2 1 1000000
.ends 0603_744761220A_200n
*******
.subckt 0603_744761220GA_200n 1 2
C1 1 N7 96.5504f
L1 1 N1 185n
L2 N1 N2 7.0859n
L3 N2 N3 4.0485n
L4 N3 N4 19.1761n
L5 N4 N5 97.5419p
L6 N5 N6 82.1736p
R1 2 N1 9.9312
R2 2 N2 6.1986
R3 2 N3 2.8562
R4 2 N4 3.5033
R5 2 N5 3.501
R6 2 N6 3.5
R7 2 N7 41.8699
R8 2 1 1000000
.ends 0603_744761220GA_200n
*******
.subckt 0603_744761221A_210n 1 2
C1 1 N7 102.9818f
L1 1 N1 190n
L2 N1 N2 8.4483n
L3 N2 N3 8.2277n
L4 N3 N4 38.8113n
L5 N4 N5 98.4496p
L6 N5 N6 82.4272p
R1 2 N1 11.1368
R2 2 N2 5.8653
R3 2 N3 4.2003
R4 2 N4 3.9309
R5 2 N5 3.927
R6 2 N6 3.9254
R7 2 N7 44.8088
R8 2 1 1000000
.ends 0603_744761221A_210n
*******
.subckt 0603_744761221GA_210n 1 2
C1 1 N7 102.9818f
L1 1 N1 190n
L2 N1 N2 8.4483n
L3 N2 N3 8.2277n
L4 N3 N4 38.8113n
L5 N4 N5 98.4496p
L6 N5 N6 82.4272p
R1 2 N1 11.1368
R2 2 N2 5.8653
R3 2 N3 4.2003
R4 2 N4 3.9309
R5 2 N5 3.927
R6 2 N6 3.9254
R7 2 N7 44.8088
R8 2 1 1000000
.ends 0603_744761221GA_210n
*******
.subckt 0603_744761222A_220n 1 2
C1 1 N7 80.2203f
L1 1 N1 200n
L2 N1 N2 7.0382n
L3 N2 N3 7.8692n
L4 N3 N4 38.8470n
L5 N4 N5 98.4794p
L6 N5 N6 82.4613p
R1 2 N1 11.1293
R2 2 N2 5.854
R3 2 N3 4.1963
R4 2 N4 3.933
R5 2 N5 3.9291
R6 2 N6 3.9275
R7 2 N7 44.6968
R8 2 1 1000000
.ends 0603_744761222A_220n
*******
.subckt 0603_744761222GA_220n 1 2
C1 1 N7 80.2203f
L1 1 N1 200n
L2 N1 N2 7.0382n
L3 N2 N3 7.8692n
L4 N3 N4 38.8470n
L5 N4 N5 98.4794p
L6 N5 N6 82.4613p
R1 2 N1 11.1293
R2 2 N2 5.854
R3 2 N3 4.1963
R4 2 N4 3.933
R5 2 N5 3.9291
R6 2 N6 3.9275
R7 2 N7 44.6968
R8 2 1 1000000
.ends 0603_744761222GA_220n
*******
.subckt 0603_744761224A_240n 1 2
C1 1 N7 94.7374f
L1 1 N1 215n
L2 N1 N2 8.1578n
L3 N2 N3 5.5993n
L4 N3 N4 38.9348n
L5 N4 N5 98.4708p
L6 N5 N6 82.4470p
R1 2 N1 11.1678
R2 2 N2 5.8063
R3 2 N3 4.1342
R4 2 N4 3.9497
R5 2 N5 3.9458
R6 2 N6 3.9442
R7 2 N7 44.8679
R8 2 1 1000000
.ends 0603_744761224A_240n
*******
.subckt 0603_744761224GA_240n 1 2
C1 1 N7 94.7374f
L1 1 N1 215n
L2 N1 N2 8.1578n
L3 N2 N3 5.5993n
L4 N3 N4 38.9348n
L5 N4 N5 98.4708p
L6 N5 N6 82.4470p
R1 2 N1 11.1678
R2 2 N2 5.8063
R3 2 N3 4.1342
R4 2 N4 3.9497
R5 2 N5 3.9458
R6 2 N6 3.9442
R7 2 N7 44.8679
R8 2 1 1000000
.ends 0603_744761224GA_240n
*******
.subckt 0603_744761227A_270n 1 2
C1 1 N7 75.3613f
L1 1 N1 245n
L2 N1 N2 10.5897n
L3 N2 N3 2.0424n
L4 N3 N4 53.1169n
L5 N4 N5 102.4122p
L6 N5 N6 86.5553p
R1 2 N1 13.1232
R2 2 N2 5.9777
R3 2 N3 5.2399
R4 2 N4 4.4028
R5 2 N5 4.3982
R6 2 N6 4.3963
R7 2 N7 49.253
R8 2 1 1000000
.ends 0603_744761227A_270n
*******
.subckt 0603_744761227GA_270n 1 2
C1 1 N7 75.3613f
L1 1 N1 245n
L2 N1 N2 10.5897n
L3 N2 N3 2.0424n
L4 N3 N4 53.1169n
L5 N4 N5 102.4122p
L6 N5 N6 86.5553p
R1 2 N1 13.1232
R2 2 N2 5.9777
R3 2 N3 5.2399
R4 2 N4 4.4028
R5 2 N5 4.3982
R6 2 N6 4.3963
R7 2 N7 49.253
R8 2 1 1000000
.ends 0603_744761227GA_270n
*******
.subckt 0603_744761233A_330n 1 2
C1 1 N7 0.3p
L1 1 N1 300n
L2 N1 N2 3.7096n
L3 N2 N3 3.9081n
L4 N3 N4 25.0400n
L5 N4 N5 180.4856p
L6 N5 N6 113.5229p
R1 2 N1 18.9649
R2 2 N2 43.3125
R3 2 N3 9.5356
R4 2 N4 6.6161
R5 2 N5 6.5169
R6 2 N6 6.4737
R7 2 N7 155.5859
R8 2 1 1000000
.ends 0603_744761233A_330n
*******
.subckt 0603_744761233GA_330n 1 2
C1 1 N7 0.3p
L1 1 N1 300n
L2 N1 N2 3.7096n
L3 N2 N3 3.9081n
L4 N3 N4 25.0400n
L5 N4 N5 180.4856p
L6 N5 N6 113.5229p
R1 2 N1 18.9649
R2 2 N2 43.3125
R3 2 N3 9.5356
R4 2 N4 6.6161
R5 2 N5 6.5169
R6 2 N6 6.4737
R7 2 N7 155.5859
R8 2 1 1000000
.ends 0603_744761233GA_330n
*******
.subckt 0603_744761239A_390n 1 2
C1 1 N7 308.8089f
L1 1 N1 360n
L2 N1 N2 21.5077n
L3 N2 N3 9.1105n
L4 N3 N4 42.3740n
L5 N4 N5 183.5558p
L6 N5 N6 117.4379p
R1 2 N1 19.6527
R2 2 N2 5.3675
R3 2 N3 9.5915
R4 2 N4 6.6284
R5 2 N5 6.5295
R6 2 N6 6.4865
R7 2 N7 25.865
R8 2 1 1000000
.ends 0603_744761239A_390n
*******
.subckt 0603_744761239GA_390n 1 2
C1 1 N7 308.8089f
L1 1 N1 360n
L2 N1 N2 21.5077n
L3 N2 N3 9.1105n
L4 N3 N4 42.3740n
L5 N4 N5 183.5558p
L6 N5 N6 117.4379p
R1 2 N1 19.6527
R2 2 N2 5.3675
R3 2 N3 9.5915
R4 2 N4 6.6284
R5 2 N5 6.5295
R6 2 N6 6.4865
R7 2 N7 25.865
R8 2 1 1000000
.ends 0603_744761239GA_390n
*******
.subckt 0603_744761247A_470n 1 2
C1 1 N7 88.6450f
L1 1 N1 440n
L2 N1 N2 11.2420n
L3 N2 N3 5.8068n
L4 N3 N4 34.9792n
L5 N4 N5 1.0010n
L6 N5 N6 1.0007n
R1 2 N1 46.4339
R2 2 N2 25.1672
R3 2 N3 13.657
R4 2 N4 13.4098
R5 2 N5 9.5927
R6 2 N6 8.5608
R7 2 N7 49.154
R8 2 1 10g
.ends 0603_744761247A_470n
*******
.subckt 0603_744761256A_560n 1 2
C1 1 N7 448.4260f
L1 1 N1 520n
L2 N1 N2 14.1825n
L3 N2 N3 31.7466n
L4 N3 N4 18.8024n
L5 N4 N5 1.0006n
L6 N5 N6 1.0008n
R1 2 N1 46.8669
R2 2 N2 26.5125
R3 2 N3 11.6335
R4 2 N4 11.0512
R5 2 N5 9.5526
R6 2 N6 8.5104
R7 2 N7 51.4228
R8 2 1 10g
.ends 0603_744761256A_560n
*******
.subckt 0603_744761268A_680n 1 2
C1 1 N7 188.5298f
L1 1 N1 600n
L2 N1 N2 36.9371n
L3 N2 N3 37.1922n
L4 N3 N4 58.2271n
L5 N4 N5 201.8001p
L6 N5 N6 144.1100p
R1 2 N1 39.4757
R2 2 N2 9.1957
R3 2 N3 9.7351
R4 2 N4 6.8518
R5 2 N5 6.7595
R6 2 N6 6.7194
R7 2 N7 37.6872
R8 2 1 1000000
.ends 0603_744761268A_680n
*******
.subckt 0603_744761282A_820n 1 2
C1 1 N7 479.2933f
L1 1 N1 770n
L2 N1 N2 19.1190n
L3 N2 N3 64.1035n
L4 N3 N4 30.7245n
L5 N4 N5 1.0015n
L6 N5 N6 1.0018n
R1 2 N1 49.2693
R2 2 N2 32.9437
R3 2 N3 7.8632
R4 2 N4 6.1563
R5 2 N5 9.5041
R6 2 N6 8.449
R7 2 N7 53.3258
R8 2 1 10g
.ends 0603_744761282A_820n
*******
.subckt 0603_744761310A_1000n 1 2
C1 1 N7 159.5551f
L1 1 N1 850n
L2 N1 N2 39.2620n
L3 N2 N3 59.0386n
L4 N3 N4 595.0270n
L5 N4 N5 1.4585n
L6 N5 N6 759.7885p
R1 2 N1 145.1307
R2 2 N2 32.9239
R3 2 N3 5.8618
R4 2 N4 6.6698
R5 2 N5 6.5722
R6 2 N6 6.5297
R7 2 N7 216.8879
R8 2 1 1000000
.ends 0603_744761310A_1000n
*******
.subckt 0805_744760022A_2.2n 1 2
C1 1 N7 283.0942f
L1 1 N1 2.1n
L2 N1 N2 61.5732p
L3 N2 N3 39.0918p
L4 N3 N4 102.4450p
L5 N4 N5 76.1894p
L6 N5 N6 53.8139p
R1 2 N1 394.4571m
R2 2 N2 471.3327m
R3 2 N3 101.7490m
R4 2 N4 138.1444m
R5 2 N5 94.4479m
R6 2 N6 86.4002m
R7 2 N7 1.9436
R8 2 1 1000000
.ends 0805_744760022A_2.2n
*******
.subckt 0805_744760027A_2.7n 1 2
C1 1 N7 265.8269f
L1 1 N1 2.6n
L2 N1 N2 112.8250p
L3 N2 N3 94.2236p
L4 N3 N4 124.0286p
L5 N4 N5 89.3975p
L6 N5 N6 57.0326p
R1 2 N1 709.1234m
R2 2 N2 618.1986m
R3 2 N3 140.4318m
R4 2 N4 454.1599m
R5 2 N5 103.8070m
R6 2 N6 93.5764m
R7 2 N7 1.9251
R8 2 1 1000000
.ends 0805_744760027A_2.7n
*******
.subckt 0805_744760033A_3.3n 1 2
C1 1 N7 181.7100f
L1 1 N1 3.2n
L2 N1 N2 48.3167p
L3 N2 N3 94.5939p
L4 N3 N4 145.6333p
L5 N4 N5 89.5607p
L6 N5 N6 57.0748p
R1 2 N1 684.1296m
R2 2 N2 615.9728m
R3 2 N3 171.7416m
R4 2 N4 455.7370m
R5 2 N5 116.7713m
R6 2 N6 93.6959m
R7 2 N7 1.9245
R8 2 1 1000000
.ends 0805_744760033A_3.3n
*******
.subckt 0805_744760039A_3.9n 1 2
C1 1 N7 111.8813f
L1 1 N1 3.7n
L2 N1 N2 90.1937p
L3 N2 N3 96.8643p
L4 N3 N4 322.0827p
L5 N4 N5 91.0418p
L6 N5 N6 57.6865p
R1 2 N1 653.9486m
R2 2 N2 620.6902m
R3 2 N3 317.5129m
R4 2 N4 475.0603m
R5 2 N5 227.1312m
R6 2 N6 96.1644m
R7 2 N7 1.9228
R8 2 1 1000000
.ends 0805_744760039A_3.9n
*******
.subckt 0805_744760047A_4.7n 1 2
C1 1 N7 146.9545f
L1 1 N1 4.5n
L2 N1 N2 99.6252p
L3 N2 N3 98.3439p
L4 N3 N4 573.3935p
L5 N4 N5 93.6332p
L6 N5 N6 59.2500p
R1 2 N1 612.1612m
R2 2 N2 601.2706m
R3 2 N3 270.6141m
R4 2 N4 526.7901m
R5 2 N5 418.6338m
R6 2 N6 105.9778m
R7 2 N7 1.9245
R8 2 1 1000000
.ends 0805_744760047A_4.7n
*******
.subckt 0805_744760051A_5.1n 1 2
C1 1 N7 169.5947f
L1 1 N1 4.8n
L2 N1 N2 147.7174p
L3 N2 N3 97.7174p
L4 N3 N4 561.3136p
L5 N4 N5 93.5571p
L6 N5 N6 59.2069p
R1 2 N1 667.2044m
R2 2 N2 593.0803m
R3 2 N3 218.5749m
R4 2 N4 525.5863m
R5 2 N5 417.6868m
R6 2 N6 105.8825m
R7 2 N7 1.9246
R8 2 1 1000000
.ends 0805_744760051A_5.1n
*******
.subckt 0805_744760056A_5.6n 1 2
C1 1 N7 180.8470f
L1 1 N1 5.3n
L2 N1 N2 161.0627p
L3 N2 N3 97.2181p
L4 N3 N4 557.6864p
L5 N4 N5 93.5329p
L6 N5 N6 59.1935p
R1 2 N1 742.9475m
R2 2 N2 587.8807m
R3 2 N3 212.6290m
R4 2 N4 525.8044m
R5 2 N5 418.3081m
R6 2 N6 105.9943m
R7 2 N7 1.9245
R8 2 1 1000000
.ends 0805_744760056A_5.6n
*******
.subckt 0805_744760056GA_5.6n 1 2
C1 1 N7 180.8470f
L1 1 N1 5.3n
L2 N1 N2 161.0627p
L3 N2 N3 97.2181p
L4 N3 N4 557.6864p
L5 N4 N5 93.5329p
L6 N5 N6 59.1935p
R1 2 N1 742.9475m
R2 2 N2 587.8807m
R3 2 N3 212.6290m
R4 2 N4 525.8044m
R5 2 N5 418.3081m
R6 2 N6 105.9943m
R7 2 N7 1.9245
R8 2 1 1000000
.ends 0805_744760056GA_5.6n
*******
.subckt 0805_744760068A_6.8n 1 2
C1 1 N7 119.7699f
L1 1 N1 6.5n
L2 N1 N2 122.1756p
L3 N2 N3 100.3315p
L4 N3 N4 625.4600p
L5 N4 N5 93.9679p
L6 N5 N6 59.4557p
R1 2 N1 665.3988m
R2 2 N2 641.0144m
R3 2 N3 498.5459m
R4 2 N4 535.5975m
R5 2 N5 428.6163m
R6 2 N6 107.2947m
R7 2 N7 1.9232
R8 2 1 1000000
.ends 0805_744760068A_6.8n
*******
.subckt 0805_744760068GA_6.8n 1 2
C1 1 N7 119.7699f
L1 1 N1 6.5n
L2 N1 N2 122.1756p
L3 N2 N3 100.3315p
L4 N3 N4 625.4600p
L5 N4 N5 93.9679p
L6 N5 N6 59.4557p
R1 2 N1 665.3988m
R2 2 N2 641.0144m
R3 2 N3 498.5459m
R4 2 N4 535.5975m
R5 2 N5 428.6163m
R6 2 N6 107.2947m
R7 2 N7 1.9232
R8 2 1 1000000
.ends 0805_744760068GA_6.8n
*******
.subckt 0805_744760082A_8.2n 1 2
C1 1 N7 185.1580f
L1 1 N1 7.85n
L2 N1 N2 217.8462p
L3 N2 N3 99.8149p
L4 N3 N4 630.0985p
L5 N4 N5 94.0522p
L6 N5 N6 59.5242p
R1 2 N1 796.7458m
R2 2 N2 622.9716m
R3 2 N3 467.7717m
R4 2 N4 539.1143m
R5 2 N5 434.2692m
R6 2 N6 108.1412m
R7 2 N7 1.9249
R8 2 1 1000000
.ends 0805_744760082A_8.2n
*******
.subckt 0805_744760082GA_8.2n 1 2
C1 1 N7 185.1580f
L1 1 N1 7.85n
L2 N1 N2 217.8462p
L3 N2 N3 99.8149p
L4 N3 N4 630.0985p
L5 N4 N5 94.0522p
L6 N5 N6 59.5242p
R1 2 N1 796.7458m
R2 2 N2 622.9716m
R3 2 N3 467.7717m
R4 2 N4 539.1143m
R5 2 N5 434.2692m
R6 2 N6 108.1412m
R7 2 N7 1.9249
R8 2 1 1000000
.ends 0805_744760082GA_8.2n
*******
.subckt 0805_744760110A_10n 1 2
C1 1 N7 219.4880f
L1 1 N1 9.7n
L2 N1 N2 289.7404p
L3 N2 N3 100.0542p
L4 N3 N4 661.5486p
L5 N4 N5 94.2936p
L6 N5 N6 59.6842p
R1 2 N1 886.4651m
R2 2 N2 633.4141m
R3 2 N3 486.7748m
R4 2 N4 545.4587m
R5 2 N5 441.9917m
R6 2 N6 109.2160m
R7 2 N7 1.9294
R8 2 1 1000000
.ends 0805_744760110A_10n
*******
.subckt 0805_744760110GA_10n 1 2
C1 1 N7 219.4880f
L1 1 N1 9.7n
L2 N1 N2 289.7404p
L3 N2 N3 100.0542p
L4 N3 N4 661.5486p
L5 N4 N5 94.2936p
L6 N5 N6 59.6842p
R1 2 N1 886.4651m
R2 2 N2 633.4141m
R3 2 N3 486.7748m
R4 2 N4 545.4587m
R5 2 N5 441.9917m
R6 2 N6 109.2160m
R7 2 N7 1.9294
R8 2 1 1000000
.ends 0805_744760110GA_10n
*******
.subckt 0805_744760112A_12n 1 2
C1 1 N7 153.3229f
L1 1 N1 11.7n
L2 N1 N2 407.3100p
L3 N2 N3 103.0651p
L4 N3 N4 935.1684p
L5 N4 N5 96.3045p
L6 N5 N6 60.9851p
R1 2 N1 929.0744m
R2 2 N2 743.7999m
R3 2 N3 670.2271m
R4 2 N4 599.6610m
R5 2 N5 505.2864m
R6 2 N6 118.6342m
R7 2 N7 1.9388
R8 2 1 1000000
.ends 0805_744760112A_12n
*******
.subckt 0805_744760112GA_12n 1 2
C1 1 N7 153.3229f
L1 1 N1 11.7n
L2 N1 N2 407.3100p
L3 N2 N3 103.0651p
L4 N3 N4 935.1684p
L5 N4 N5 96.3045p
L6 N5 N6 60.9851p
R1 2 N1 929.0744m
R2 2 N2 743.7999m
R3 2 N3 670.2271m
R4 2 N4 599.6610m
R5 2 N5 505.2864m
R6 2 N6 118.6342m
R7 2 N7 1.9388
R8 2 1 1000000
.ends 0805_744760112GA_12n
*******
.subckt 0805_744760115A_15n 1 2
C1 1 N7 205.2469f
L1 1 N1 14.6n
L2 N1 N2 457.9816p
L3 N2 N3 103.2962p
L4 N3 N4 1.0260n
L5 N4 N5 97.0138p
L6 N5 N6 61.4578p
R1 2 N1 1.266
R2 2 N2 748.4897m
R3 2 N3 687.0761m
R4 2 N4 621.9851m
R5 2 N5 531.7582m
R6 2 N6 123.0240m
R7 2 N7 1.9768
R8 2 1 1000000
.ends 0805_744760115A_15n
*******
.subckt 0805_744760115GA_15n 1 2
C1 1 N7 205.2469f
L1 1 N1 14.6n
L2 N1 N2 457.9816p
L3 N2 N3 103.2962p
L4 N3 N4 1.0260n
L5 N4 N5 97.0138p
L6 N5 N6 61.4578p
R1 2 N1 1.266
R2 2 N2 748.4897m
R3 2 N3 687.0761m
R4 2 N4 621.9851m
R5 2 N5 531.7582m
R6 2 N6 123.0240m
R7 2 N7 1.9768
R8 2 1 1000000
.ends 0805_744760115GA_15n
*******
.subckt 0805_744760118A_18n 1 2
C1 1 N7 133.7155f
L1 1 N1 17.6n
L2 N1 N2 345.4904p
L3 N2 N3 103.0207p
L4 N3 N4 1.0245n
L5 N4 N5 97.0080p
L6 N5 N6 61.4541p
R1 2 N1 1.2276
R2 2 N2 734.2501m
R3 2 N3 678.1061m
R4 2 N4 622.0457m
R5 2 N5 531.9886m
R6 2 N6 123.0753m
R7 2 N7 1.9767
R8 2 1 1000000
.ends 0805_744760118A_18n
*******
.subckt 0805_744760118GA_18n 1 2
C1 1 N7 133.7155f
L1 1 N1 17.6n
L2 N1 N2 345.4904p
L3 N2 N3 103.0207p
L4 N3 N4 1.0245n
L5 N4 N5 97.0080p
L6 N5 N6 61.4541p
R1 2 N1 1.2276
R2 2 N2 734.2501m
R3 2 N3 678.1061m
R4 2 N4 622.0457m
R5 2 N5 531.9886m
R6 2 N6 123.0753m
R7 2 N7 1.9767
R8 2 1 1000000
.ends 0805_744760118GA_18n
*******
.subckt 0805_744760122A_22n 1 2
C1 1 N7 125.6488f
L1 1 N1 21n
L2 N1 N2 905.8708p
L3 N2 N3 106.9745p
L4 N3 N4 1.2229n
L5 N4 N5 98.9922p
L6 N5 N6 62.7572p
R1 2 N1 1.3296
R2 2 N2 903.5546m
R3 2 N3 857.6462m
R4 2 N4 681.4068m
R5 2 N5 598.1705m
R6 2 N6 134.4052m
R7 2 N7 2.0007
R8 2 1 1000000
.ends 0805_744760122A_22n
*******
.subckt 0805_744760122GA_22n 1 2
C1 1 N7 125.6488f
L1 1 N1 21n
L2 N1 N2 905.8708p
L3 N2 N3 106.9745p
L4 N3 N4 1.2229n
L5 N4 N5 98.9922p
L6 N5 N6 62.7572p
R1 2 N1 1.3296
R2 2 N2 903.5546m
R3 2 N3 857.6462m
R4 2 N4 681.4068m
R5 2 N5 598.1705m
R6 2 N6 134.4052m
R7 2 N7 2.0007
R8 2 1 1000000
.ends 0805_744760122GA_22n
*******
.subckt 0805_744760127A_27n 1 2
C1 1 N7 176.5700f
L1 1 N1 26.2n
L2 N1 N2 776.2439p
L3 N2 N3 110.0620p
L4 N3 N4 1.2229n
L5 N4 N5 102.8478p
L6 N5 N6 65.3543p
R1 2 N1 1.7176
R2 2 N2 981.7006m
R3 2 N3 984.1757m
R4 2 N4 794.4310m
R5 2 N5 719.7253m
R6 2 N6 156.8785m
R7 2 N7 2.0855
R8 2 1 1000000
.ends 0805_744760127A_27n
*******
.subckt 0805_744760127GA_27n 1 2
C1 1 N7 176.5700f
L1 1 N1 26.2n
L2 N1 N2 776.2439p
L3 N2 N3 110.0620p
L4 N3 N4 1.2229n
L5 N4 N5 102.8478p
L6 N5 N6 65.3543p
R1 2 N1 1.7176
R2 2 N2 981.7006m
R3 2 N3 984.1757m
R4 2 N4 794.4310m
R5 2 N5 719.7253m
R6 2 N6 156.8785m
R7 2 N7 2.0855
R8 2 1 1000000
.ends 0805_744760127GA_27n
*******
.subckt 0805_744760133A_33n 1 2
C1 1 N7 179.1460f
L1 1 N1 32n
L2 N1 N2 1.1088n
L3 N2 N3 145.3441p
R1 2 N1 2.08
R2 2 N2 1.8125
R3 2 N3 1.4013
R7 2 N7 2.1814
R8 2 1 1000000
.ends 0805_744760133A_33n
*******
.subckt 0805_744760133GA_33n 1 2
C1 1 N7 179.1460f
L1 1 N1 32n
L2 N1 N2 1.1088n
L3 N2 N3 145.3441p
R1 2 N1 2.08
R2 2 N2 1.8125
R3 2 N3 1.4013
R7 2 N7 2.1814
R8 2 1 1000000
.ends 0805_744760133GA_33n
*******
.subckt 0805_744760136A_36n 1 2
C1 1 N7 145.4401f
L1 1 N1 35.5n
L2 N1 N2 1.1127n
L3 N2 N3 145.4552p
R1 2 N1 2.2457
R2 2 N2 1.7999
R3 2 N3 1.3896
R7 2 N7 2.2222
R8 2 1 1000000
.ends 0805_744760136A_36n
*******
.subckt 0805_744760136GA_36n 1 2
C1 1 N7 145.4401f
L1 1 N1 35.5n
L2 N1 N2 1.1127n
L3 N2 N3 145.4552p
R1 2 N1 2.2457
R2 2 N2 1.7999
R3 2 N3 1.3896
R7 2 N7 2.2222
R8 2 1 1000000
.ends 0805_744760136GA_36n
*******
.subckt 0805_744760139A_39n 1 2
C1 1 N7 131.2261f
L1 1 N1 37n
L2 N1 N2 768.4217p
L3 N2 N3 18.7678p
L4 N3 N4 1.4486n
L5 N4 N5 20.2786p
L6 N5 N6 100.2641p
R1 2 N1 2.8546
R2 2 N2 4.8233
R3 2 N3 2.9263
R4 2 N4 878.9766m
R5 2 N5 828.1977m
R6 2 N6 726.8619m
R7 2 N7 3.5313
R8 2 1 1000000
.ends 0805_744760139A_39n
*******
.subckt 0805_744760139GA_39n 1 2
C1 1 N7 131.2261f
L1 1 N1 37n
L2 N1 N2 768.4217p
L3 N2 N3 18.7678p
L4 N3 N4 1.4486n
L5 N4 N5 20.2786p
L6 N5 N6 100.2641p
R1 2 N1 2.8546
R2 2 N2 4.8233
R3 2 N3 2.9263
R4 2 N4 878.9766m
R5 2 N5 828.1977m
R6 2 N6 726.8619m
R7 2 N7 3.5313
R8 2 1 1000000
.ends 0805_744760139GA_39n
*******
.subckt 0805_744760143A_43n 1 2
C1 1 N7 142.3480f
L1 1 N1 38n
L2 N1 N2 918.7399p
L3 N2 N3 207.5538p
L4 N3 N4 11.9580n
L5 N4 N5 97.2603p
L6 N5 N6 65.2641p
R1 2 N1 2.8048
R2 2 N2 4.9331
R3 2 N3 3.1926
R4 2 N4 817.9804m
R5 2 N5 743.6095m
R6 2 N6 576.9804m
R7 2 N7 3.515
R8 2 1 1000000
.ends 0805_744760143A_43n
*******
.subckt 0805_744760143GA_43n 1 2
C1 1 N7 142.3480f
L1 1 N1 38n
L2 N1 N2 918.7399p
L3 N2 N3 207.5538p
L4 N3 N4 11.9580n
L5 N4 N5 97.2603p
L6 N5 N6 65.2641p
R1 2 N1 2.8048
R2 2 N2 4.9331
R3 2 N3 3.1926
R4 2 N4 817.9804m
R5 2 N5 743.6095m
R6 2 N6 576.9804m
R7 2 N7 3.515
R8 2 1 1000000
.ends 0805_744760143GA_43n
*******
.subckt 0805_744760147A_47n 1 2
C1 1 N7 176.8813f
L1 1 N1 43n
L2 N1 N2 894.7222p
L3 N2 N3 188.0372p
L4 N3 N4 1.9822n
L5 N4 N5 13.5482p
L6 N5 N6 64.4546p
R1 2 N1 2.647
R2 2 N2 4.6132
R3 2 N3 2.3618
R4 2 N4 785.5399m
R5 2 N5 709.9673m
R6 2 N6 530.6681m
R7 2 N7 2.0904
R8 2 1 1000000
.ends 0805_744760147A_47n
*******
.subckt 0805_744760147GA_47n 1 2
C1 1 N7 176.8813f
L1 1 N1 43n
L2 N1 N2 894.7222p
L3 N2 N3 188.0372p
L4 N3 N4 1.9822n
L5 N4 N5 13.5482p
L6 N5 N6 64.4546p
R1 2 N1 2.647
R2 2 N2 4.6132
R3 2 N3 2.3618
R4 2 N4 785.5399m
R5 2 N5 709.9673m
R6 2 N6 530.6681m
R7 2 N7 2.0904
R8 2 1 1000000
.ends 0805_744760147GA_47n
*******
.subckt 0805_744760156A_56n 1 2
C1 1 N7 137.4379f
L1 1 N1 52n
L2 N1 N2 2.0026n
L3 N2 N3 174.3144p
L4 N3 N4 7.0919n
L5 N4 N5 14.0722p
L6 N5 N6 64.6026p
R1 2 N1 2.9976
R2 2 N2 4.6032
R3 2 N3 2.3236
R4 2 N4 870.0859m
R5 2 N5 810.2154m
R6 2 N6 687.3630m
R7 2 N7 2.1529
R8 2 1 1000000
.ends 0805_744760156A_56n
*******
.subckt 0805_744760156GA_56n 1 2
C1 1 N7 137.4379f
L1 1 N1 52n
L2 N1 N2 2.0026n
L3 N2 N3 174.3144p
L4 N3 N4 7.0919n
L5 N4 N5 14.0722p
L6 N5 N6 64.6026p
R1 2 N1 2.9976
R2 2 N2 4.6032
R3 2 N3 2.3236
R4 2 N4 870.0859m
R5 2 N5 810.2154m
R6 2 N6 687.3630m
R7 2 N7 2.1529
R8 2 1 1000000
.ends 0805_744760156GA_56n
*******
.subckt 0805_744760168A_68n 1 2
C1 1 N7 145.4642f
L1 1 N1 62n
L2 N1 N2 1.8534n
L3 N2 N3 161.1445p
L4 N3 N4 3.7068n
L5 N4 N5 14.0369p
L6 N5 N6 64.5747p
R1 2 N1 2.9818
R2 2 N2 4.5978
R3 2 N3 2.3003
R4 2 N4 828.8488m
R5 2 N5 762.1436m
R6 2 N6 617.6620m
R7 2 N7 2.1009
R8 2 1 1000000
.ends 0805_744760168A_68n
*******
.subckt 0805_744760168GA_68n 1 2
C1 1 N7 145.4642f
L1 1 N1 62n
L2 N1 N2 1.8534n
L3 N2 N3 161.1445p
L4 N3 N4 3.7068n
L5 N4 N5 14.0369p
L6 N5 N6 64.5747p
R1 2 N1 2.9818
R2 2 N2 4.5978
R3 2 N3 2.3003
R4 2 N4 828.8488m
R5 2 N5 762.1436m
R6 2 N6 617.6620m
R7 2 N7 2.1009
R8 2 1 1000000
.ends 0805_744760168GA_68n
*******
.subckt 0805_744760182A_82n 1 2
C1 1 N7 143.9062f
L1 1 N1 75n
L2 N1 N2 3.3238n
L3 N2 N3 188.6327p
L4 N3 N4 10.0191n
L5 N4 N5 14.3819p
L6 N5 N6 64.6747p
R1 2 N1 3.5491
R2 2 N2 4.5991
R3 2 N3 2.3086
R4 2 N4 952.0781m
R5 2 N5 903.6480m
R6 2 N6 812.8171m
R7 2 N7 2.1611
R8 2 1 1000000
.ends 0805_744760182A_82n
*******
.subckt 0805_744760182GA_82n 1 2
C1 1 N7 143.9062f
L1 1 N1 75n
L2 N1 N2 3.3238n
L3 N2 N3 188.6327p
L4 N3 N4 10.0191n
L5 N4 N5 14.3819p
L6 N5 N6 64.6747p
R1 2 N1 3.5491
R2 2 N2 4.5991
R3 2 N3 2.3086
R4 2 N4 952.0781m
R5 2 N5 903.6480m
R6 2 N6 812.8171m
R7 2 N7 2.1611
R8 2 1 1000000
.ends 0805_744760182GA_82n
*******
.subckt 0805_744760191A_91n 1 2
C1 1 N7 138.6745f
L1 1 N1 83n
L2 N1 N2 3.9189n
L3 N2 N3 193.1871p
L4 N3 N4 10.9843n
L5 N4 N5 14.5328p
L6 N5 N6 64.7108p
R1 2 N1 3.7443
R2 2 N2 4.6005
R3 2 N3 2.3142
R4 2 N4 977.8751m
R5 2 N5 932.1083m
R6 2 N6 847.4702m
R7 2 N7 2.1839
R8 2 1 1000000
.ends 0805_744760191A_91n
*******
.subckt 0805_744760191GA_91n 1 2
C1 1 N7 138.6745f
L1 1 N1 83n
L2 N1 N2 3.9189n
L3 N2 N3 193.1871p
L4 N3 N4 10.9843n
L5 N4 N5 14.5328p
L6 N5 N6 64.7108p
R1 2 N1 3.7443
R2 2 N2 4.6005
R3 2 N3 2.3142
R4 2 N4 977.8751m
R5 2 N5 932.1083m
R6 2 N6 847.4702m
R7 2 N7 2.1839
R8 2 1 1000000
.ends 0805_744760191GA_91n
*******
.subckt 0805_744760210A_100n 1 2
C1 1 N7 193.6123f
L1 1 N1 90n
L2 N1 N2 3.6981n
L3 N2 N3 185.1060p
L4 N3 N4 10.8857n
L5 N4 N5 14.5237p
L6 N5 N6 64.7087p
R1 2 N1 3.908
R2 2 N2 4.5952
R3 2 N3 2.2931
R4 2 N4 983.0668m
R5 2 N5 937.8266m
R6 2 N6 854.3977m
R7 2 N7 2.2116
R8 2 1 1000000
.ends 0805_744760210A_100n
*******
.subckt 0805_744760210GA_100n 1 2
C1 1 N7 193.6123f
L1 1 N1 90n
L2 N1 N2 3.6981n
L3 N2 N3 185.1060p
L4 N3 N4 10.8857n
L5 N4 N5 14.5237p
L6 N5 N6 64.7087p
R1 2 N1 3.908
R2 2 N2 4.5952
R3 2 N3 2.2931
R4 2 N4 983.0668m
R5 2 N5 937.8266m
R6 2 N6 854.3977m
R7 2 N7 2.2116
R8 2 1 1000000
.ends 0805_744760210GA_100n
*******
.subckt 0805_744760212A_120n 1 2
C1 1 N7 172.4332f
L1 1 N1 110n
L2 N1 N2 4.5578n
L3 N2 N3 178.1949p
L4 N3 N4 11.0643n
L5 N4 N5 15.1803p
L6 N5 N6 64.8576p
R1 2 N1 4.3259
R2 2 N2 4.5782
R3 2 N3 2.2212
R4 2 N4 1.0367
R5 2 N5 996.3688m
R6 2 N6 923.9227m
R7 2 N7 2.224
R8 2 1 1000000
.ends 0805_744760212A_120n
*******
.subckt 0805_744760212GA_120n 1 2
C1 1 N7 172.4332f
L1 1 N1 110n
L2 N1 N2 4.5578n
L3 N2 N3 178.1949p
L4 N3 N4 11.0643n
L5 N4 N5 15.1803p
L6 N5 N6 64.8576p
R1 2 N1 4.3259
R2 2 N2 4.5782
R3 2 N3 2.2212
R4 2 N4 1.0367
R5 2 N5 996.3688m
R6 2 N6 923.9227m
R7 2 N7 2.224
R8 2 1 1000000
.ends 0805_744760212GA_120n
*******
.subckt 0805_744760215A_150n 1 2
C1 1 N7 177.3022f
L1 1 N1 135n
L2 N1 N2 5.8282n
L3 N2 N3 187.8851p
L4 N3 N4 12.4729n
L5 N4 N5 16.5430p
L6 N5 N6 65.1815p
R1 2 N1 4.9215
R2 2 N2 4.5701
R3 2 N3 2.1845
R4 2 N4 1.1154
R5 2 N5 1.081
R6 2 N6 1.0209
R7 2 N7 2.2739
R8 2 1 1000000
.ends 0805_744760215A_150n
*******
.subckt 0805_744760215GA_150n 1 2
C1 1 N7 177.3022f
L1 1 N1 135n
L2 N1 N2 5.8282n
L3 N2 N3 187.8851p
L4 N3 N4 12.4729n
L5 N4 N5 16.5430p
L6 N5 N6 65.1815p
R1 2 N1 4.9215
R2 2 N2 4.5701
R3 2 N3 2.1845
R4 2 N4 1.1154
R5 2 N5 1.081
R6 2 N6 1.0209
R7 2 N7 2.2739
R8 2 1 1000000
.ends 0805_744760215GA_150n
*******
.subckt 0805_744760218A_180n 1 2
C1 1 N7 172.8852f
L1 1 N1 165n
L2 N1 N2 7.8777n
L3 N2 N3 221.1119p
L4 N3 N4 15.7816n
L5 N4 N5 19.1152p
L6 N5 N6 65.8579p
R1 2 N1 5.8378
R2 2 N2 4.575
R3 2 N3 2.2039
R4 2 N4 1.253
R5 2 N5 1.2261
R6 2 N6 1.1806
R7 2 N7 2.3707
R8 2 1 1000000
.ends 0805_744760218A_180n
*******
.subckt 0805_744760218GA_180n 1 2
C1 1 N7 172.8852f
L1 1 N1 165n
L2 N1 N2 7.8777n
L3 N2 N3 221.1119p
L4 N3 N4 15.7816n
L5 N4 N5 19.1152p
L6 N5 N6 65.8579p
R1 2 N1 5.8378
R2 2 N2 4.575
R3 2 N3 2.2039
R4 2 N4 1.253
R5 2 N5 1.2261
R6 2 N6 1.1806
R7 2 N7 2.3707
R8 2 1 1000000
.ends 0805_744760218GA_180n
*******
.subckt 0805_744760222A_220n 1 2
C1 1 N7 60.3568f
L1 1 N1 210n
L2 N1 N2 6.6378n
L3 N2 N3 522.8939p
L4 N3 N4 17.8667n
L5 N4 N5 101.1970p
L6 N5 N6 66.5250p
R1 2 N1 14.962
R2 2 N2 5.8415
R3 2 N3 5.2294
R4 2 N4 4.4029
R5 2 N5 4.3984
R6 2 N6 4.3965
R7 2 N7 49.29
R8 2 1 1000000
.ends 0805_744760222A_220n
*******
.subckt 0805_744760222GA_220n 1 2
C1 1 N7 60.3568f
L1 1 N1 210n
L2 N1 N2 6.6378n
L3 N2 N3 522.8939p
L4 N3 N4 17.8667n
L5 N4 N5 101.1970p
L6 N5 N6 66.5250p
R1 2 N1 14.962
R2 2 N2 5.8415
R3 2 N3 5.2294
R4 2 N4 4.4029
R5 2 N5 4.3984
R6 2 N6 4.3965
R7 2 N7 49.29
R8 2 1 1000000
.ends 0805_744760222GA_220n
*******
.subckt 0805_744760227A_270n 1 2
C1 1 N7 65.9663f
L1 1 N1 250n
L2 N1 N2 8.5809n
L3 N2 N3 471.8863p
L4 N3 N4 23.7013n
L5 N4 N5 101.4607p
L6 N5 N6 66.5256p
R1 2 N1 15.068
R2 2 N2 5.8402
R3 2 N3 5.2279
R4 2 N4 4.403
R5 2 N5 4.3985
R6 2 N6 4.3966
R7 2 N7 49.2889
R8 2 1 1000000
.ends 0805_744760227A_270n
*******
.subckt 0805_744760227GA_270n 1 2
C1 1 N7 65.9663f
L1 1 N1 250n
L2 N1 N2 8.5809n
L3 N2 N3 471.8863p
L4 N3 N4 23.7013n
L5 N4 N5 101.4607p
L6 N5 N6 66.5256p
R1 2 N1 15.068
R2 2 N2 5.8402
R3 2 N3 5.2279
R4 2 N4 4.403
R5 2 N5 4.3985
R6 2 N6 4.3966
R7 2 N7 49.2889
R8 2 1 1000000
.ends 0805_744760227GA_270n
*******
.subckt 0805_744760233A_330n 1 2
C1 1 N7 83.3061f
L1 1 N1 310n
L2 N1 N2 12.8190n
L3 N2 N3 759.5331p
L4 N3 N4 35.4501n
L5 N4 N5 101.9993p
L6 N5 N6 66.5271p
R1 2 N1 14.7696
R2 2 N2 5.846
R3 2 N3 5.2351
R4 2 N4 4.4046
R5 2 N5 4.4001
R6 2 N6 4.3982
R7 2 N7 49.2925
R8 2 1 1000000
.ends 0805_744760233A_330n
*******
.subckt 0805_744760233GA_330n 1 2
C1 1 N7 83.3061f
L1 1 N1 310n
L2 N1 N2 12.8190n
L3 N2 N3 759.5331p
L4 N3 N4 35.4501n
L5 N4 N5 101.9993p
L6 N5 N6 66.5271p
R1 2 N1 14.7696
R2 2 N2 5.846
R3 2 N3 5.2351
R4 2 N4 4.4046
R5 2 N5 4.4001
R6 2 N6 4.3982
R7 2 N7 49.2925
R8 2 1 1000000
.ends 0805_744760233GA_330n
*******
.subckt 0805_744760239A_390n 1 2
C1 1 N7 138.6278f
L1 1 N1 365n
L2 N1 N2 9.9330n
L3 N2 N3 2.0379n
L4 N3 N4 24.2012n
L5 N4 N5 31.5293p
L6 N5 N6 69.3148p
R1 2 N1 15.0525
R2 2 N2 12.9906
R3 2 N3 12.2367
R4 2 N4 5.0885
R5 2 N5 5.0948
R6 2 N6 5.1064
R7 2 N7 3.5112
R8 2 1 1000000
.ends 0805_744760239A_390n
*******
.subckt 0805_744760239GA_390n 1 2
C1 1 N7 138.6278f
L1 1 N1 365n
L2 N1 N2 9.9330n
L3 N2 N3 2.0379n
L4 N3 N4 24.2012n
L5 N4 N5 31.5293p
L6 N5 N6 69.3148p
R1 2 N1 15.0525
R2 2 N2 12.9906
R3 2 N3 12.2367
R4 2 N4 5.0885
R5 2 N5 5.0948
R6 2 N6 5.1064
R7 2 N7 3.5112
R8 2 1 1000000
.ends 0805_744760239GA_390n
*******
.subckt 0805_7447602470A_470n 1 2
C1 1 N7 300.6151f
L1 1 N1 440n
L2 N1 N2 18.2484n
L3 N2 N3 7.4881n
L4 N3 N4 46.5226n
L5 N4 N5 1.0022n
L6 N5 N6 1.0022n
R1 2 N1 49.1505
R2 2 N2 32.2514
R3 2 N3 7.4442
R4 2 N4 2.0109
R5 2 N5 9.4949
R6 2 N6 8.4374
R7 2 N7 55.2898
R8 2 1 10g
.ends 0805_7447602470A_470n
*******
.subckt 0805_7447602560A_560n 1 2
C1 1 N7 158.6203f
L1 1 N1 530n
L2 N1 N2 18.4815n
L3 N2 N3 15.7345n
L4 N3 N4 67.3500n
L5 N4 N5 1.0027n
L6 N5 N6 1.0025n
R1 2 N1 49.1872
R2 2 N2 32.2832
R3 2 N3 8.7525
R4 2 N4 3.6958
R5 2 N5 9.4964
R6 2 N6 8.4392
R7 2 N7 55.7968
R8 2 1 10g
.ends 0805_7447602560A_560n
*******
.subckt 0805_7447602620A_620n 1 2
C1 1 N7 374.7521f
L1 1 N1 580n
L2 N1 N2 18.5875n
L3 N2 N3 21.6723n
L4 N3 N4 69.8015n
L5 N4 N5 1.0026n
L6 N5 N6 1.0023n
R1 2 N1 49.2018
R2 2 N2 32.3273
R3 2 N3 8.859
R4 2 N4 3.8426
R5 2 N5 9.4966
R6 2 N6 8.4395
R7 2 N7 55.8259
R8 2 1 10g
.ends 0805_7447602620A_620n
*******
.subckt 0805_7447602680A_680n 1 2
C1 1 N7 299.9001f
L1 1 N1 640n
L2 N1 N2 18.6377n
L3 N2 N3 27.2681n
L4 N3 N4 67.6580n
L5 N4 N5 1.0027n
L6 N5 N6 1.0024n
R1 2 N1 49.1914
R2 2 N2 32.3246
R3 2 N3 8.8938
R4 2 N4 3.6851
R5 2 N5 9.4964
R6 2 N6 8.4392
R7 2 N7 55.8063
R8 2 1 10g
.ends 0805_7447602680A_680n
*******
.subckt 0805_7447602820A_820n 1 2
C1 1 N7 392.3243f
L1 1 N1 780n
L2 N1 N2 18.9312n
L3 N2 N3 41.9285n
L4 N3 N4 57.3860n
L5 N4 N5 1.0025n
L6 N5 N6 1.0024n
R1 2 N1 49.2521
R2 2 N2 32.5078
R3 2 N3 8.8827
R4 2 N4 2.83
R5 2 N5 9.4953
R6 2 N6 8.4378
R7 2 N7 55.8726
R8 2 1 10g
.ends 0805_7447602820A_820n
*******
.subckt 0805_7447603100A_1000n 1 2
C1 1 N7 321.3970f
L1 1 N1 970n
L2 N1 N2 26.2072n
L3 N2 N3 59.5963n
L4 N3 N4 37.9513n
L5 N4 N5 1.0055n
L6 N5 N6 1.0058n
R1 2 N1 54.2392
R2 2 N2 42.0066
R3 2 N3 13.1987
R4 2 N4 16.2089
R5 2 N5 9.6181
R6 2 N6 8.5926
R7 2 N7 57.8314
R8 2 1 10g
.ends 0805_7447603100A_1000n
*******
.subckt 0805_7447603120A_1200n 1 2
C1 1 N7 386.7332f
L1 1 N1 1160n
L2 N1 N2 31.1907n
L3 N2 N3 79.8927n
L4 N3 N4 40.4710n
L5 N4 N5 1.0084n
L6 N5 N6 1.0082n
R1 2 N1 58.6432
R2 2 N2 48.5362
R3 2 N3 18.732
R4 2 N4 20.536
R5 2 N5 9.7507
R6 2 N6 8.7581
R7 2 N7 59.5493
R8 2 1 10g
.ends 0805_7447603120A_1200n
*******
.subckt 0805_7447603150A_1500n 1 2
C1 1 N7 261.5429f
L1 1 N1 1400n
L2 N1 N2 48.3637n
L3 N2 N3 31.9729n
L4 N3 N4 70.2203n
L5 N4 N5 1.0293n
L6 N5 N6 1.0243n
R1 2 N1 74.768
R2 2 N2 65.4601
R3 2 N3 38.0258
R4 2 N4 44.7014
R5 2 N5 11.847
R6 2 N6 11.2268
R7 2 N7 69.7816
R8 2 1 10g
.ends 0805_7447603150A_1500n
*******
.subckt 0805_7447603180A_1800n 1 2
C1 1 N7 254.8407f
L1 1 N1 1650n
L2 N1 N2 51.1609n
L3 N2 N3 61.4284n
L4 N3 N4 59.4592n
L5 N4 N5 1.0367n
L6 N5 N6 1.0316n
R1 2 N1 77.2754
R2 2 N2 67.8266
R3 2 N3 40.9591
R4 2 N4 47.1026
R5 2 N5 12.1931
R6 2 N6 11.6106
R7 2 N7 71.9328
R8 2 1 10g
.ends 0805_7447603180A_1800n
*******
.subckt 1008_744762033A_3.3n 1 2
C1 1 N7 258.8890f
L1 1 N1 3.2n
L2 N1 N2 74.6295p
L3 N2 N3 27.5037p
L4 N3 N4 178.7950p
L5 N4 N5 125.8937p
L6 N5 N6 64.4396p
R1 2 N1 496.4370m
R2 2 N2 652.0149m
R3 2 N3 174.5643m
R4 2 N4 196.4350m
R5 2 N5 175.6405m
R6 2 N6 166.1640m
R7 2 N7 2.0868
R8 2 1 1000000
.ends 1008_744762033A_3.3n
*******
.subckt 1008_744762039A_3.9n 1 2
C1 1 N7 307.3090f
L1 1 N1 3.8n
L2 N1 N2 171.8081p
L3 N2 N3 64.6854p
L4 N3 N4 227.3111p
L5 N4 N5 150.1826p
L6 N5 N6 64.5035p
R1 2 N1 613.4031m
R2 2 N2 647.3909m
R3 2 N3 222.0463m
R4 2 N4 225.6419m
R5 2 N5 195.1920m
R6 2 N6 183.4104m
R7 2 N7 2.0882
R8 2 1 1000000
.ends 1008_744762039A_3.9n
*******
.subckt 1008_744762068A_6.8n 1 2
C1 1 N7 154.0665f
L1 1 N1 6.7n
L2 N1 N2 166.2730p
L3 N2 N3 108.7064p
L4 N3 N4 318.1466p
L5 N4 N5 191.3683p
L6 N5 N6 64.6221p
R1 2 N1 661.4449m
R2 2 N2 648.3710m
R3 2 N3 309.3671m
R4 2 N4 273.2139m
R5 2 N5 225.5854m
R6 2 N6 211.0042m
R7 2 N7 2.0817
R8 2 1 1000000
.ends 1008_744762068A_6.8n
*******
.subckt 1008_744762068GA_6.8n 1 2
C1 1 N7 154.0665f
L1 1 N1 6.7n
L2 N1 N2 166.2730p
L3 N2 N3 108.7064p
L4 N3 N4 318.1466p
L5 N4 N5 191.3683p
L6 N5 N6 64.6221p
R1 2 N1 661.4449m
R2 2 N2 648.3710m
R3 2 N3 309.3671m
R4 2 N4 273.2139m
R5 2 N5 225.5854m
R6 2 N6 211.0042m
R7 2 N7 2.0817
R8 2 1 1000000
.ends 1008_744762068GA_6.8n
*******
.subckt 1008_744762082A_8.2n 1 2
C1 1 N7 134.7654f
L1 1 N1 8.1n
L2 N1 N2 189.4028p
L3 N2 N3 181.8662p
L4 N3 N4 408.3459p
L5 N4 N5 308.8976p
L6 N5 N6 66.4859p
R1 2 N1 762.2513m
R2 2 N2 418.0814m
R3 2 N3 232.8557m
R4 2 N4 313.9906m
R5 2 N5 846.3900m
R6 2 N6 552.8978m
R7 2 N7 3.4553
R8 2 1 1000000
.ends 1008_744762082A_8.2n
*******
.subckt 1008_744762082GA_8.2n 1 2
C1 1 N7 134.7654f
L1 1 N1 8.1n
L2 N1 N2 189.4028p
L3 N2 N3 181.8662p
L4 N3 N4 408.3459p
L5 N4 N5 308.8976p
L6 N5 N6 66.4859p
R1 2 N1 762.2513m
R2 2 N2 418.0814m
R3 2 N3 232.8557m
R4 2 N4 313.9906m
R5 2 N5 846.3900m
R6 2 N6 552.8978m
R7 2 N7 3.4553
R8 2 1 1000000
.ends 1008_744762082GA_8.2n
*******
.subckt 1008_744762110A_10n 1 2
C1 1 N7 181.1045f
L1 1 N1 9.5n
L2 N1 N2 359.5564p
L3 N2 N3 233.2733p
L4 N3 N4 427.9970p
L5 N4 N5 312.9171p
L6 N5 N6 66.5085p
R1 2 N1 878.4726m
R2 2 N2 448.4753m
R3 2 N3 292.8569m
R4 2 N4 322.8625m
R5 2 N5 846.4481m
R6 2 N6 552.6441m
R7 2 N7 3.4561
R8 2 1 1000000
.ends 1008_744762110A_10n
*******
.subckt 1008_744762110GA_10n 1 2
C1 1 N7 181.1045f
L1 1 N1 9.5n
L2 N1 N2 359.5564p
L3 N2 N3 233.2733p
L4 N3 N4 427.9970p
L5 N4 N5 312.9171p
L6 N5 N6 66.5085p
R1 2 N1 878.4726m
R2 2 N2 448.4753m
R3 2 N3 292.8569m
R4 2 N4 322.8625m
R5 2 N5 846.4481m
R6 2 N6 552.6441m
R7 2 N7 3.4561
R8 2 1 1000000
.ends 1008_744762110GA_10n
*******
.subckt 1008_744762112A_12n 1 2
C1 1 N7 146.8195f
L1 1 N1 11.5n
L2 N1 N2 277.8637p
L3 N2 N3 275.2129p
L4 N3 N4 445.2785p
L5 N4 N5 316.7401p
L6 N5 N6 66.5175p
R1 2 N1 859.4485m
R2 2 N2 457.5956m
R3 2 N3 328.8614m
R4 2 N4 329.4138m
R5 2 N5 846.1378m
R6 2 N6 551.7080m
R7 2 N7 3.4563
R8 2 1 1000000
.ends 1008_744762112A_12n
*******
.subckt 1008_744762112GA_12n 1 2
C1 1 N7 146.8195f
L1 1 N1 11.5n
L2 N1 N2 277.8637p
L3 N2 N3 275.2129p
L4 N3 N4 445.2785p
L5 N4 N5 316.7401p
L6 N5 N6 66.5175p
R1 2 N1 859.4485m
R2 2 N2 457.5956m
R3 2 N3 328.8614m
R4 2 N4 329.4138m
R5 2 N5 846.1378m
R6 2 N6 551.7080m
R7 2 N7 3.4563
R8 2 1 1000000
.ends 1008_744762112GA_12n
*******
.subckt 1008_744762115A_15n 1 2
C1 1 N7 157.0687f
L1 1 N1 14.5n
L2 N1 N2 271.9509p
L3 N2 N3 303.1149p
L4 N3 N4 444.2736p
L5 N4 N5 317.1278p
L6 N5 N6 66.5239p
R1 2 N1 815.7379m
R2 2 N2 471.7354m
R3 2 N3 313.7702m
R4 2 N4 317.8127m
R5 2 N5 844.4898m
R6 2 N6 547.6468m
R7 2 N7 3.4563
R8 2 1 1000000
.ends 1008_744762115A_15n
*******
.subckt 1008_744762115GA_15n 1 2
C1 1 N7 157.0687f
L1 1 N1 14.5n
L2 N1 N2 271.9509p
L3 N2 N3 303.1149p
L4 N3 N4 444.2736p
L5 N4 N5 317.1278p
L6 N5 N6 66.5239p
R1 2 N1 815.7379m
R2 2 N2 471.7354m
R3 2 N3 313.7702m
R4 2 N4 317.8127m
R5 2 N5 844.4898m
R6 2 N6 547.6468m
R7 2 N7 3.4563
R8 2 1 1000000
.ends 1008_744762115GA_15n
*******
.subckt 1008_744762118A_18n 1 2
C1 1 N7 225.1780f
L1 1 N1 17.5n
L2 N1 N2 497.7966p
L3 N2 N3 349.6621p
L4 N3 N4 471.4224p
L5 N4 N5 322.9627p
L6 N5 N6 66.5450p
R1 2 N1 990.3641m
R2 2 N2 501.8900m
R3 2 N3 351.0477m
R4 2 N4 318.2605m
R5 2 N5 842.7047m
R6 2 N6 542.8637m
R7 2 N7 3.4575
R8 2 1 1000000
.ends 1008_744762118A_18n
*******
.subckt 1008_744762118GA_18n 1 2
C1 1 N7 225.1780f
L1 1 N1 17.5n
L2 N1 N2 497.7966p
L3 N2 N3 349.6621p
L4 N3 N4 471.4224p
L5 N4 N5 322.9627p
L6 N5 N6 66.5450p
R1 2 N1 990.3641m
R2 2 N2 501.8900m
R3 2 N3 351.0477m
R4 2 N4 318.2605m
R5 2 N5 842.7047m
R6 2 N6 542.8637m
R7 2 N7 3.4575
R8 2 1 1000000
.ends 1008_744762118GA_18n
*******
.subckt 1008_744762122A_22n 1 2
C1 1 N7 153.5785f
L1 1 N1 21n
L2 N1 N2 401.9102p
L3 N2 N3 347.0378p
L4 N3 N4 477.3577p
L5 N4 N5 324.4792p
L6 N5 N6 66.5542p
R1 2 N1 928.4318m
R2 2 N2 480.0546m
R3 2 N3 350.6736m
R4 2 N4 313.2296m
R5 2 N5 841.5736m
R6 2 N6 539.9744m
R7 2 N7 3.4565
R8 2 1 1000000
.ends 1008_744762122A_22n
*******
.subckt 1008_744762122GA_22n 1 2
C1 1 N7 153.5785f
L1 1 N1 21n
L2 N1 N2 401.9102p
L3 N2 N3 347.0378p
L4 N3 N4 477.3577p
L5 N4 N5 324.4792p
L6 N5 N6 66.5542p
R1 2 N1 928.4318m
R2 2 N2 480.0546m
R3 2 N3 350.6736m
R4 2 N4 313.2296m
R5 2 N5 841.5736m
R6 2 N6 539.9744m
R7 2 N7 3.4565
R8 2 1 1000000
.ends 1008_744762122GA_22n
*******
.subckt 1008_744762127A_27n 1 2
C1 1 N7 235.3466f
L1 1 N1 26n
L2 N1 N2 760.5796p
L3 N2 N3 1.0152n
L4 N3 N4 896.3806p
L5 N4 N5 455.4809p
L6 N5 N6 67.0501p
R1 2 N1 1.3469
R2 2 N2 856.8490m
R3 2 N3 953.0422m
R4 2 N4 762.4712m
R5 2 N5 929.8044m
R6 2 N6 717.7057m
R7 2 N7 3.4968
R8 2 1 1000000
.ends 1008_744762127A_27n
*******
.subckt 1008_744762127GA_27n 1 2
C1 1 N7 235.3466f
L1 1 N1 26n
L2 N1 N2 760.5796p
L3 N2 N3 1.0152n
L4 N3 N4 896.3806p
L5 N4 N5 455.4809p
L6 N5 N6 67.0501p
R1 2 N1 1.3469
R2 2 N2 856.8490m
R3 2 N3 953.0422m
R4 2 N4 762.4712m
R5 2 N5 929.8044m
R6 2 N6 717.7057m
R7 2 N7 3.4968
R8 2 1 1000000
.ends 1008_744762127GA_27n
*******
.subckt 1008_744762133A_33n 1 2
C1 1 N7 168.6910f
L1 1 N1 31.5n
L2 N1 N2 677.8936p
L3 N2 N3 802.4968p
L4 N3 N4 804.0651p
L5 N4 N5 423.3038p
L6 N5 N6 66.9467p
R1 2 N1 1.2068
R2 2 N2 308.2071m
R3 2 N3 798.8010m
R4 2 N4 647.1974m
R5 2 N5 873.2351m
R6 2 N6 618.7997m
R7 2 N7 3.5004
R8 2 1 1000000
.ends 1008_744762133A_33n
*******
.subckt 1008_744762133GA_33n 1 2
C1 1 N7 168.6910f
L1 1 N1 31.5n
L2 N1 N2 677.8936p
L3 N2 N3 802.4968p
L4 N3 N4 804.0651p
L5 N4 N5 423.3038p
L6 N5 N6 66.9467p
R1 2 N1 1.2068
R2 2 N2 308.2071m
R3 2 N3 798.8010m
R4 2 N4 647.1974m
R5 2 N5 873.2351m
R6 2 N6 618.7997m
R7 2 N7 3.5004
R8 2 1 1000000
.ends 1008_744762133GA_33n
*******
.subckt 1008_744762139A_39n 1 2
C1 1 N7 203.2740f
L1 1 N1 38n
L2 N1 N2 1.5622n
L3 N2 N3 1.9110n
L4 N3 N4 1.4779n
L5 N4 N5 697.7198p
L6 N5 N6 68.2205p
R1 2 N1 1.726
R2 2 N2 1.7074
R3 2 N3 1.5914
R4 2 N4 1.267
R5 2 N5 1.1436
R6 2 N6 1.0926
R7 2 N7 3.5849
R8 2 1 1000000
.ends 1008_744762139A_39n
*******
.subckt 1008_744762139GA_39n 1 2
C1 1 N7 203.2740f
L1 1 N1 38n
L2 N1 N2 1.5622n
L3 N2 N3 1.9110n
L4 N3 N4 1.4779n
L5 N4 N5 697.7198p
L6 N5 N6 68.2205p
R1 2 N1 1.726
R2 2 N2 1.7074
R3 2 N3 1.5914
R4 2 N4 1.267
R5 2 N5 1.1436
R6 2 N6 1.0926
R7 2 N7 3.5849
R8 2 1 1000000
.ends 1008_744762139GA_39n
*******
.subckt 1008_744762147A_47n 1 2
C1 1 N7 187.1203f
L1 1 N1 46n
L2 N1 N2 1.2911n
L3 N2 N3 1.9110n
L4 N3 N4 1.5623n
L5 N4 N5 740.2101p
L6 N5 N6 68.3322p
R1 2 N1 2.0169
R2 2 N2 1.5313
R3 2 N3 1.6598
R4 2 N4 1.3405
R5 2 N5 1.209
R6 2 N6 1.1626
R7 2 N7 3.6683
R8 2 1 1000000
.ends 1008_744762147A_47n
*******
.subckt 1008_744762147GA_47n 1 2
C1 1 N7 187.1203f
L1 1 N1 46n
L2 N1 N2 1.2911n
L3 N2 N3 1.9110n
L4 N3 N4 1.5623n
L5 N4 N5 740.2101p
L6 N5 N6 68.3322p
R1 2 N1 2.0169
R2 2 N2 1.5313
R3 2 N3 1.6598
R4 2 N4 1.3405
R5 2 N5 1.209
R6 2 N6 1.1626
R7 2 N7 3.6683
R8 2 1 1000000
.ends 1008_744762147GA_47n
*******
.subckt 1008_744762156A_56n 1 2
C1 1 N7 257.2154f
L1 1 N1 54n
L2 N1 N2 1.2136n
L3 N2 N3 2.1376n
L4 N3 N4 347.2515p
L5 N4 N5 721.8134p
L6 N5 N6 68.2728p
R1 2 N1 2.3751
R2 2 N2 477.1832m
R3 2 N3 1.5003
R4 2 N4 1.1955
R5 2 N5 1.0402
R6 2 N6 977.8847m
R7 2 N7 4.9999
R8 2 1 1000000
.ends 1008_744762156A_56n
*******
.subckt 1008_744762156GA_56n 1 2
C1 1 N7 257.2154f
L1 1 N1 54n
L2 N1 N2 1.2136n
L3 N2 N3 2.1376n
L4 N3 N4 347.2515p
L5 N4 N5 721.8134p
L6 N5 N6 68.2728p
R1 2 N1 2.3751
R2 2 N2 477.1832m
R3 2 N3 1.5003
R4 2 N4 1.1955
R5 2 N5 1.0402
R6 2 N6 977.8847m
R7 2 N7 4.9999
R8 2 1 1000000
.ends 1008_744762156GA_56n
*******
.subckt 1008_744762168A_68n 1 2
C1 1 N7 193.0510f
L1 1 N1 65n
L2 N1 N2 1.3983n
L3 N2 N3 1.5992n
L4 N3 N4 1.5233n
L5 N4 N5 730.6600p
L6 N5 N6 68.3061p
R1 2 N1 2.4167
R2 2 N2 603.5214m
R3 2 N3 1.5436
R4 2 N4 1.2687
R5 2 N5 1.1294
R6 2 N6 1.0764
R7 2 N7 3.9404
R8 2 1 1000000
.ends 1008_744762168A_68n
*******
.subckt 1008_744762168GA_68n 1 2
C1 1 N7 193.0510f
L1 1 N1 65n
L2 N1 N2 1.3983n
L3 N2 N3 1.5992n
L4 N3 N4 1.5233n
L5 N4 N5 730.6600p
L6 N5 N6 68.3061p
R1 2 N1 2.4167
R2 2 N2 603.5214m
R3 2 N3 1.5436
R4 2 N4 1.2687
R5 2 N5 1.1294
R6 2 N6 1.0764
R7 2 N7 3.9404
R8 2 1 1000000
.ends 1008_744762168GA_68n
*******
.subckt 1008_744762182A_82n 1 2
C1 1 N7 148.9036f
L1 1 N1 80n
L2 N1 N2 1.5838n
L3 N2 N3 1.6561n
L4 N3 N4 1.5487n
L5 N4 N5 1.5487n
L6 N5 N6 68.3935p
R1 2 N1 3.4312
R2 2 N2 820.5022m
R3 2 N3 1.4873
R4 2 N4 1.1492
R5 2 N5 964.4580m
R6 2 N6 890.8371m
R7 2 N7 4.3017
R8 2 1 1000000
.ends 1008_744762182A_82n
*******
.subckt 1008_744762182GA_82n 1 2
C1 1 N7 148.9036f
L1 1 N1 80n
L2 N1 N2 1.5838n
L3 N2 N3 1.6561n
L4 N3 N4 1.5487n
L5 N4 N5 1.5487n
L6 N5 N6 68.3935p
R1 2 N1 3.4312
R2 2 N2 820.5022m
R3 2 N3 1.4873
R4 2 N4 1.1492
R5 2 N5 964.4580m
R6 2 N6 890.8371m
R7 2 N7 4.3017
R8 2 1 1000000
.ends 1008_744762182GA_82n
*******
.subckt 1008_744762210A_100n 1 2
C1 1 N7 160.6109f
L1 1 N1 95n
L2 N1 N2 1.9043n
L3 N2 N3 1.1914n
L4 N3 N4 2.7207n
L5 N4 N5 3.0832n
L6 N5 N6 2.0638n
R1 2 N1 5.5161
R2 2 N2 4.8896
R3 2 N3 2.9794
R4 2 N4 2.7578
R5 2 N5 2.2546
R6 2 N6 2.2396
R7 2 N7 7.7857
R8 2 1 1000000
.ends 1008_744762210A_100n
*******
.subckt 1008_744762210GA_100n 1 2
C1 1 N7 160.6109f
L1 1 N1 95n
L2 N1 N2 1.9043n
L3 N2 N3 1.1914n
L4 N3 N4 2.7207n
L5 N4 N5 3.0832n
L6 N5 N6 2.0638n
R1 2 N1 5.5161
R2 2 N2 4.8896
R3 2 N3 2.9794
R4 2 N4 2.7578
R5 2 N5 2.2546
R6 2 N6 2.2396
R7 2 N7 7.7857
R8 2 1 1000000
.ends 1008_744762210GA_100n
*******
.subckt 1008_744762212A_120n 1 2
C1 1 N7 180.5203f
L1 1 N1 110n
L2 N1 N2 1.9916n
L3 N2 N3 171.8219p
L4 N3 N4 1.6406n
L5 N4 N5 2.6544n
L6 N5 N6 1.9729n
R1 2 N1 5.5201
R2 2 N2 4.8873
R3 2 N3 2.9697
R4 2 N4 2.7508
R5 2 N5 2.2512
R6 2 N6 2.2379
R7 2 N7 7.7857
R8 2 1 1000000
.ends 1008_744762212A_120n
*******
.subckt 1008_744762212GA_120n 1 2
C1 1 N7 180.5203f
L1 1 N1 110n
L2 N1 N2 1.9916n
L3 N2 N3 171.8219p
L4 N3 N4 1.6406n
L5 N4 N5 2.6544n
L6 N5 N6 1.9729n
R1 2 N1 5.5201
R2 2 N2 4.8873
R3 2 N3 2.9697
R4 2 N4 2.7508
R5 2 N5 2.2512
R6 2 N6 2.2379
R7 2 N7 7.7857
R8 2 1 1000000
.ends 1008_744762212GA_120n
*******
.subckt 1008_744762215A_150n 1 2
C1 1 N7 209.3657f
L1 1 N1 140n
L2 N1 N2 3.5326n
L3 N2 N3 177.3744p
L4 N3 N4 3.3242n
L5 N4 N5 3.2593n
L6 N5 N6 2.0910n
R1 2 N1 5.5226
R2 2 N2 4.8969
R3 2 N3 2.9961
R4 2 N4 2.7695
R5 2 N5 2.2673
R6 2 N6 2.2518
R7 2 N7 7.7854
R8 2 1 1000000
.ends 1008_744762215A_150n
*******
.subckt 1008_744762215GA_150n 1 2
C1 1 N7 209.3657f
L1 1 N1 140n
L2 N1 N2 3.5326n
L3 N2 N3 177.3744p
L4 N3 N4 3.3242n
L5 N4 N5 3.2593n
L6 N5 N6 2.0910n
R1 2 N1 5.5226
R2 2 N2 4.8969
R3 2 N3 2.9961
R4 2 N4 2.7695
R5 2 N5 2.2673
R6 2 N6 2.2518
R7 2 N7 7.7854
R8 2 1 1000000
.ends 1008_744762215GA_150n
*******
.subckt 1008_744762218A_180n 1 2
C1 1 N7 193.1000f
L1 1 N1 172n
L2 N1 N2 4.5246n
L3 N2 N3 181.0740p
L4 N3 N4 4.4839n
L5 N4 N5 3.5882n
L6 N5 N6 2.1583n
R1 2 N1 5.5047
R2 2 N2 4.9108
R3 2 N3 3.0335
R4 2 N4 2.7942
R5 2 N5 2.2962
R6 2 N6 2.2798
R7 2 N7 17.7817
R8 2 1 1000000
.ends 1008_744762218A_180n
*******
.subckt 1008_744762218GA_180n 1 2
C1 1 N7 193.1000f
L1 1 N1 172n
L2 N1 N2 4.5246n
L3 N2 N3 181.0740p
L4 N3 N4 4.4839n
L5 N4 N5 3.5882n
L6 N5 N6 2.1583n
R1 2 N1 5.5047
R2 2 N2 4.9108
R3 2 N3 3.0335
R4 2 N4 2.7942
R5 2 N5 2.2962
R6 2 N6 2.2798
R7 2 N7 17.7817
R8 2 1 1000000
.ends 1008_744762218GA_180n
*******
.subckt 1008_744762222A_220n 1 2
C1 1 N7 156.8026f
L1 1 N1 210n
L2 N1 N2 4.7562n
L3 N2 N3 1.9220n
L4 N3 N4 8.6154n
L5 N4 N5 5.2009n
L6 N5 N6 4.2055n
R1 2 N1 8.6651
R2 2 N2 4.9153
R3 2 N3 3.0695
R4 2 N4 2.8166
R5 2 N5 2.3232
R6 2 N6 2.306
R7 2 N7 27.7798
R8 2 1 1000000
.ends 1008_744762222A_220n
*******
.subckt 1008_744762222GA_220n 1 2
C1 1 N7 156.8026f
L1 1 N1 210n
L2 N1 N2 4.7562n
L3 N2 N3 1.9220n
L4 N3 N4 8.6154n
L5 N4 N5 5.2009n
L6 N5 N6 4.2055n
R1 2 N1 8.6651
R2 2 N2 4.9153
R3 2 N3 3.0695
R4 2 N4 2.8166
R5 2 N5 2.3232
R6 2 N6 2.306
R7 2 N7 27.7798
R8 2 1 1000000
.ends 1008_744762222GA_220n
*******
.subckt 1008_744762227A_270n 1 2
C1 1 N7 134.9807f
L1 1 N1 255n
L2 N1 N2 5.9174n
L3 N2 N3 2.4737n
L4 N3 N4 8.6718n
L5 N4 N5 5.2147n
L6 N5 N6 4.2084n
R1 2 N1 8.6661
R2 2 N2 4.9196
R3 2 N3 3.0743
R4 2 N4 2.8176
R5 2 N5 2.3241
R6 2 N6 2.3068
R7 2 N7 27.7796
R8 2 1 1000000
.ends 1008_744762227A_270n
*******
.subckt 1008_744762227GA_270n 1 2
C1 1 N7 134.9807f
L1 1 N1 255n
L2 N1 N2 5.9174n
L3 N2 N3 2.4737n
L4 N3 N4 8.6718n
L5 N4 N5 5.2147n
L6 N5 N6 4.2084n
R1 2 N1 8.6661
R2 2 N2 4.9196
R3 2 N3 3.0743
R4 2 N4 2.8176
R5 2 N5 2.3241
R6 2 N6 2.3068
R7 2 N7 27.7796
R8 2 1 1000000
.ends 1008_744762227GA_270n
*******
.subckt 1008_744762233A_330n 1 2
C1 1 N7 166.9531f
L1 1 N1 320n
L2 N1 N2 8.7552n
L3 N2 N3 4.6165n
L4 N3 N4 16.4431n
L5 N4 N5 11.1334n
L6 N5 N6 4.0890n
R1 2 N1 8.6723
R2 2 N2 4.9113
R3 2 N3 3.0421
R4 2 N4 2.8054
R5 2 N5 9.3131
R6 2 N6 7.8736
R7 2 N7 27.7777
R8 2 1 1000000
.ends 1008_744762233A_330n
*******
.subckt 1008_744762233GA_330n 1 2
C1 1 N7 166.9531f
L1 1 N1 320n
L2 N1 N2 8.7552n
L3 N2 N3 4.6165n
L4 N3 N4 16.4431n
L5 N4 N5 11.1334n
L6 N5 N6 4.0890n
R1 2 N1 8.6723
R2 2 N2 4.9113
R3 2 N3 3.0421
R4 2 N4 2.8054
R5 2 N5 9.3131
R6 2 N6 7.8736
R7 2 N7 27.7777
R8 2 1 1000000
.ends 1008_744762233GA_330n
*******
.subckt 1008_744762239A_390n 1 2
C1 1 N7 178.5846f
L1 1 N1 370n
L2 N1 N2 11.5605n
L3 N2 N3 5.4024n
L4 N3 N4 16.4967n
L5 N4 N5 11.1427n
L6 N5 N6 4.0926n
R1 2 N1 8.6862
R2 2 N2 4.9288
R3 2 N3 3.0538
R4 2 N4 2.814
R5 2 N5 9.3138
R6 2 N6 7.8746
R7 2 N7 27.7776
R8 2 1 1000000
.ends 1008_744762239A_390n
*******
.subckt 1008_744762239GA_390n 1 2
C1 1 N7 178.5846f
L1 1 N1 370n
L2 N1 N2 11.5605n
L3 N2 N3 5.4024n
L4 N3 N4 16.4967n
L5 N4 N5 11.1427n
L6 N5 N6 4.0926n
R1 2 N1 8.6862
R2 2 N2 4.9288
R3 2 N3 3.0538
R4 2 N4 2.814
R5 2 N5 9.3138
R6 2 N6 7.8746
R7 2 N7 27.7776
R8 2 1 1000000
.ends 1008_744762239GA_390n
*******
.subckt 1008_744762247A_470n 1 2
C1 1 N7 145.0718f
L1 1 N1 450n
L2 N1 N2 6.1595n
L3 N2 N3 3.1132n
L4 N3 N4 3.8323n
L5 N4 N5 10.5609n
L6 N5 N6 16.2914n
R1 2 N1 19.0285
R2 2 N2 21.5766
R3 2 N3 23.4772
R4 2 N4 11.6865
R5 2 N5 9.4736
R6 2 N6 8.0228
R7 2 N7 47.7774
R8 2 1 1000000
.ends 1008_744762247A_470n
*******
.subckt 1008_744762247GA_470n 1 2
C1 1 N7 145.0718f
L1 1 N1 450n
L2 N1 N2 6.1595n
L3 N2 N3 3.1132n
L4 N3 N4 3.8323n
L5 N4 N5 10.5609n
L6 N5 N6 16.2914n
R1 2 N1 19.0285
R2 2 N2 21.5766
R3 2 N3 23.4772
R4 2 N4 11.6865
R5 2 N5 9.4736
R6 2 N6 8.0228
R7 2 N7 47.7774
R8 2 1 1000000
.ends 1008_744762247GA_470n
*******
.subckt 1008_744762256A_560n 1 2
C1 1 N7 143.7792f
L1 1 N1 520n
L2 N1 N2 8.4301n
L3 N2 N3 4.2493n
L4 N3 N4 3.8223n
L5 N4 N5 9.6340n
L6 N5 N6 15.9713n
R1 2 N1 19.0263
R2 2 N2 21.5739
R3 2 N3 23.4772
R4 2 N4 11.665
R5 2 N5 9.4428
R6 2 N6 7.9929
R7 2 N7 47.7775
R8 2 1 1000000
.ends 1008_744762256A_560n
*******
.subckt 1008_744762256GA_560n 1 2
C1 1 N7 143.7792f
L1 1 N1 520n
L2 N1 N2 8.4301n
L3 N2 N3 4.2493n
L4 N3 N4 3.8223n
L5 N4 N5 9.6340n
L6 N5 N6 15.9713n
R1 2 N1 19.0263
R2 2 N2 21.5739
R3 2 N3 23.4772
R4 2 N4 11.665
R5 2 N5 9.4428
R6 2 N6 7.9929
R7 2 N7 47.7775
R8 2 1 1000000
.ends 1008_744762256GA_560n
*******
.subckt 1008_744762268A_680n 1 2
C1 1 N7 179.5018f
L1 1 N1 600n
L2 N1 N2 7.7623n
L3 N2 N3 7.2331n
L4 N3 N4 8.5562n
L5 N4 N5 13.3598n
L6 N5 N6 16.5293n
R1 2 N1 19.0323
R2 2 N2 21.5912
R3 2 N3 23.4825
R4 2 N4 11.7478
R5 2 N5 9.5305
R6 2 N6 8.072
R7 2 N7 47.7765
R8 2 1 1000000
.ends 1008_744762268A_680n
*******
.subckt 1008_744762268GA_680n 1 2
C1 1 N7 179.5018f
L1 1 N1 600n
L2 N1 N2 7.7623n
L3 N2 N3 7.2331n
L4 N3 N4 8.5562n
L5 N4 N5 13.3598n
L6 N5 N6 16.5293n
R1 2 N1 19.0323
R2 2 N2 21.5912
R3 2 N3 23.4825
R4 2 N4 11.7478
R5 2 N5 9.5305
R6 2 N6 8.072
R7 2 N7 47.7765
R8 2 1 1000000
.ends 1008_744762268GA_680n
*******
.subckt 1008_744762275A_750n 1 2
C1 1 N7 186.0994f
L1 1 N1 700n
L2 N1 N2 9.8413n
L3 N2 N3 11.5325n
L4 N3 N4 12.7937n
L5 N4 N5 15.2669n
L6 N5 N6 16.5975n
R1 2 N1 19.0378
R2 2 N2 21.6059
R3 2 N3 23.4879
R4 2 N4 11.7894
R5 2 N5 9.5559
R6 2 N6 8.0883
R7 2 N7 47.7753
R8 2 1 1000000
.ends 1008_744762275A_750n
*******
.subckt 1008_744762275GA_750n 1 2
C1 1 N7 186.0994f
L1 1 N1 700n
L2 N1 N2 9.8413n
L3 N2 N3 11.5325n
L4 N3 N4 12.7937n
L5 N4 N5 15.2669n
L6 N5 N6 16.5975n
R1 2 N1 19.0378
R2 2 N2 21.6059
R3 2 N3 23.4879
R4 2 N4 11.7894
R5 2 N5 9.5559
R6 2 N6 8.0883
R7 2 N7 47.7753
R8 2 1 1000000
.ends 1008_744762275GA_750n
*******
.subckt 1008_744762282A_820n 1 2
C1 1 N7 176.7473f
L1 1 N1 770n
L2 N1 N2 11.2194n
L3 N2 N3 13.7355n
L4 N3 N4 14.5850n
L5 N4 N5 15.9010n
L6 N5 N6 16.6499n
R1 2 N1 19.039
R2 2 N2 21.614
R3 2 N3 23.4916
R4 2 N4 11.8032
R5 2 N5 9.5607
R6 2 N6 8.089
R7 2 N7 47.7745
R8 2 1 1000000
.ends 1008_744762282A_820n
*******
.subckt 1008_744762282GA_820n 1 2
C1 1 N7 176.7473f
L1 1 N1 770n
L2 N1 N2 11.2194n
L3 N2 N3 13.7355n
L4 N3 N4 14.5850n
L5 N4 N5 15.9010n
L6 N5 N6 16.6499n
R1 2 N1 19.039
R2 2 N2 21.614
R3 2 N3 23.4916
R4 2 N4 11.8032
R5 2 N5 9.5607
R6 2 N6 8.089
R7 2 N7 47.7745
R8 2 1 1000000
.ends 1008_744762282GA_820n
*******
.subckt 1008_744762291A_910n 1 2
C1 1 N7 191.6803f
L1 1 N1 870n
L2 N1 N2 12.9293n
L3 N2 N3 16.7459n
L4 N3 N4 16.7803n
L5 N4 N5 16.5258n
L6 N5 N6 16.7053n
R1 2 N1 19.0403
R2 2 N2 21.6287
R3 2 N3 23.4989
R4 2 N4 11.8178
R5 2 N5 9.5625
R6 2 N6 8.0858
R7 2 N7 47.7729
R8 2 1 1000000
.ends 1008_744762291A_910n
*******
.subckt 1008_744762291GA_910n 1 2
C1 1 N7 191.6803f
L1 1 N1 870n
L2 N1 N2 12.9293n
L3 N2 N3 16.7459n
L4 N3 N4 16.7803n
L5 N4 N5 16.5258n
L6 N5 N6 16.7053n
R1 2 N1 19.0403
R2 2 N2 21.6287
R3 2 N3 23.4989
R4 2 N4 11.8178
R5 2 N5 9.5625
R6 2 N6 8.0858
R7 2 N7 47.7729
R8 2 1 1000000
.ends 1008_744762291GA_910n
*******
.subckt 1008_744762310A_1000n 1 2
C1 1 N7 188.5030f
L1 1 N1 950n
L2 N1 N2 12.9293n
L3 N2 N3 16.7460n
L4 N3 N4 16.7806n
L5 N4 N5 16.5259n
L6 N5 N6 16.7053n
R1 2 N1 19.04
R2 2 N2 21.6286
R3 2 N3 23.4989
R4 2 N4 11.8178
R5 2 N5 9.5624
R6 2 N6 8.0857
R7 2 N7 47.7729
R8 2 1 1000000
.ends 1008_744762310A_1000n
*******
.subckt 1008_744762310GA_1000n 1 2
C1 1 N7 188.5030f
L1 1 N1 950n
L2 N1 N2 12.9293n
L3 N2 N3 16.7460n
L4 N3 N4 16.7806n
L5 N4 N5 16.5259n
L6 N5 N6 16.7053n
R1 2 N1 19.04
R2 2 N2 21.6286
R3 2 N3 23.4989
R4 2 N4 11.8178
R5 2 N5 9.5624
R6 2 N6 8.0857
R7 2 N7 47.7729
R8 2 1 1000000
.ends 1008_744762310GA_1000n
*******
