**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminium Electrolyte Capacitors
* Matchcode:             WCAP-ATG5
* Library Type:          LTspice
* Version:               rev21a
* Created/modified by:   Ella
* Date and Time:         2022/11/18
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
.subckt 860020272001_22uF 1 2
Rser 1 3 1.44057897855
Lser 2 4 3.319934374E-09
C1 3 4 0.000022
Rpar 3 4 3333333.33333333
.ends 860020272001_22uF
*******
.subckt 860020272002_33uF 1 2
Rser 1 3 1.77224030686
Lser 2 4 3.460288413E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860020272002_33uF
*******
.subckt 860020272003_47uF 1 2
Rser 1 3 0.982709897838
Lser 2 4 4.140092263E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860020272003_47uF
*******
.subckt 860020272004_68uF 1 2
Rser 1 3 0.902109942493
Lser 2 4 3.47146856E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860020272004_68uF
*******
.subckt 860020272005_100uF 1 2
Rser 1 3 0.749886262101
Lser 2 4 4.173860292E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860020272005_100uF
*******
.subckt 860020272006_120uF 1 2
Rser 1 3 0.694443910842
Lser 2 4 3.658356583E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860020272006_120uF
*******
.subckt 860020272007_150uF 1 2
Rser 1 3 0.459959572682
Lser 2 4 3.764931838E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860020272007_150uF
*******
.subckt 860020273008_180uF 1 2
Rser 1 3 0.38
Lser 2 4 0.0000000188
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860020273008_180uF
*******
.subckt 860020273009_220uF 1 2
Rser 1 3 0.335
Lser 2 4 0.0000000208
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860020273009_220uF
*******
.subckt 860020273010_330uF 1 2
Rser 1 3 0.32698
Lser 2 4 8.713025952E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860020273010_330uF
*******
.subckt 860020273011_470uF 1 2
Rser 1 3 0.275
Lser 2 4 0.0000000187
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860020273011_470uF
*******
.subckt 860020274012_560uF 1 2
Rser 1 3 0.22
Lser 2 4 0.0000000289
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860020274012_560uF
*******
.subckt 860020274013_680uF 1 2
Rser 1 3 0.109
Lser 2 4 0.0000000258
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860020274013_680uF
*******
.subckt 860020274017_1.5mF 1 2
Rser 1 3 0.093
Lser 2 4 0.0000000299
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860020274017_1.5mF
*******
.subckt 860020275014_820uF 1 2
Rser 1 3 0.147
Lser 2 4 0.0000000206
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860020275014_820uF
*******
.subckt 860020275015_1mF 1 2
Rser 1 3 0.112
Lser 2 4 0.0000000228
C1 3 4 0.001
Rpar 3 4 100000
.ends 860020275015_1mF
*******
.subckt 860020275016_1.2mF 1 2
Rser 1 3 0.082
Lser 2 4 0.0000000251
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860020275016_1.2mF
*******
.subckt 860020275018_1.5mF 1 2
Rser 1 3 0.092
Lser 2 4 0.0000000262
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860020275018_1.5mF
*******
.subckt 860020275019_1.8mF 1 2
Rser 1 3 0.077
Lser 2 4 0.0000000255
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860020275019_1.8mF
*******
.subckt 860020275020_2.2mF 1 2
Rser 1 3 0.0655
Lser 2 4 0.0000000255
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860020275020_2.2mF
*******
.subckt 860020275021_2.7mF 1 2
Rser 1 3 0.0475
Lser 2 4 0.00000002434
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860020275021_2.7mF
*******
.subckt 860020278022_2.7mF 1 2
Rser 1 3 0.056
Lser 2 4 0.0000000265
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860020278022_2.7mF
*******
.subckt 860020278023_3.3mF 1 2
Rser 1 3 0.054
Lser 2 4 0.0000000259
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860020278023_3.3mF
*******
.subckt 860020278024_3.9mF 1 2
Rser 1 3 0.0455
Lser 2 4 0.0000000301
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860020278024_3.9mF
*******
.subckt 860020278025_4.7mF 1 2
Rser 1 3 0.043
Lser 2 4 0.0000000335
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860020278025_4.7mF
*******
.subckt 860020280026_5.6mF 1 2
Rser 1 3 0.033
Lser 2 4 0.000000035
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860020280026_5.6mF
*******
.subckt 860020280027_6.8mF 1 2
Rser 1 3 0.032
Lser 2 4 0.000000034
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860020280027_6.8mF
*******
.subckt 860020280028_8.2mF 1 2
Rser 1 3 0.0245
Lser 2 4 0.000000036
C1 3 4 0.0082
Rpar 3 4 12195.1219512195
.ends 860020280028_8.2mF
*******
.subckt 860020280029_10mF 1 2
Rser 1 3 0.0215
Lser 2 4 0.000000035
C1 3 4 0.01
Rpar 3 4 10000
.ends 860020280029_10mF
*******
.subckt 860020280030_12mF 1 2
Rser 1 3 0.021
Lser 2 4 0.0000000346
C1 3 4 0.012
Rpar 3 4 8333.33333333333
.ends 860020280030_12mF
*******
.subckt 860020281031_15mF 1 2
Rser 1 3 0.024
Lser 2 4 0.0000000362
C1 3 4 0.015
Rpar 3 4 6666.66666666667
.ends 860020281031_15mF
*******
.subckt 860020281032_18mF 1 2
Rser 1 3 0.02574
Lser 2 4 1.8246849327E-08
C1 3 4 0.018
Rpar 3 4 5555.55555555556
.ends 860020281032_18mF
*******
.subckt 860020372001_10uF 1 2
Rser 1 3 1.95182658193
Lser 2 4 4.159236184E-09
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 860020372001_10uF
*******
.subckt 860020372002_22uF 1 2
Rser 1 3 1.29358667564
Lser 2 4 3.756560656E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860020372002_22uF
*******
.subckt 860020372003_33uF 1 2
Rser 1 3 0.914336183608
Lser 2 4 3.799036286E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860020372003_33uF
*******
.subckt 860020372004_47uF 1 2
Rser 1 3 0.713834150585
Lser 2 4 4.196289743E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860020372004_47uF
*******
.subckt 860020372005_68uF 1 2
Rser 1 3 0.769103156896
Lser 2 4 3.629232947E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860020372005_68uF
*******
.subckt 860020372006_100uF 1 2
Rser 1 3 0.41
Lser 2 4 0.0000000162
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860020372006_100uF
*******
.subckt 860020373007_120uF 1 2
Rser 1 3 0.515044153466
Lser 2 4 4.791506411E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860020373007_120uF
*******
.subckt 860020373008_150uF 1 2
Rser 1 3 0.400204976739
Lser 2 4 4.907053114E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860020373008_150uF
*******
.subckt 860020373009_180uF 1 2
Rser 1 3 0.29
Lser 2 4 0.0000000184
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860020373009_180uF
*******
.subckt 860020373010_220uF 1 2
Rser 1 3 0.355
Lser 2 4 0.0000000173
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860020373010_220uF
*******
.subckt 860020373011_330uF 1 2
Rser 1 3 0.285
Lser 2 4 0.0000000213
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860020373011_330uF
*******
.subckt 860020374012_470uF 1 2
Rser 1 3 0.195
Lser 2 4 0.0000000197
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860020374012_470uF
*******
.subckt 860020374014_680uF 1 2
Rser 1 3 0.103
Lser 2 4 0.0000000225
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860020374014_680uF
*******
.subckt 860020375013_560uF 1 2
Rser 1 3 0.158
Lser 2 4 0.0000000227
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860020375013_560uF
*******
.subckt 860020375015_680uF 1 2
Rser 1 3 0.144
Lser 2 4 0.0000000247
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860020375015_680uF
*******
.subckt 860020375016_820uF 1 2
Rser 1 3 0.131
Lser 2 4 0.000000024
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860020375016_820uF
*******
.subckt 860020375017_1mF 1 2
Rser 1 3 0.071
Lser 2 4 0.0000000243
C1 3 4 0.001
Rpar 3 4 100000
.ends 860020375017_1mF
*******
.subckt 860020375018_1.2mF 1 2
Rser 1 3 0.077
Lser 2 4 0.0000000256
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860020375018_1.2mF
*******
.subckt 860020375019_1.5mF 1 2
Rser 1 3 0.051
Lser 2 4 0.0000000264
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860020375019_1.5mF
*******
.subckt 860020378020_1.8mF 1 2
Rser 1 3 0.063
Lser 2 4 0.0000000276
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860020378020_1.8mF
*******
.subckt 860020378021_2.2mF 1 2
Rser 1 3 0.053
Lser 2 4 0.000000019
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860020378021_2.2mF
*******
.subckt 860020378022_2.7mF 1 2
Rser 1 3 0.053
Lser 2 4 0.0000000285
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860020378022_2.7mF
*******
.subckt 860020378023_3.3mF 1 2
Rser 1 3 0.053
Lser 2 4 0.0000000258
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860020378023_3.3mF
*******
.subckt 860020380024_3.9mF 1 2
Rser 1 3 0.032
Lser 2 4 0.00000003
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860020380024_3.9mF
*******
.subckt 860020380025_4.7mF 1 2
Rser 1 3 0.0336
Lser 2 4 0.0000000234
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860020380025_4.7mF
*******
.subckt 860020380026_5.6mF 1 2
Rser 1 3 0.027
Lser 2 4 0.0000000296
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860020380026_5.6mF
*******
.subckt 860020380027_6.8mF 1 2
Rser 1 3 0.026
Lser 2 4 0.0000000358
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860020380027_6.8mF
*******
.subckt 860020380028_8.2mF 1 2
Rser 1 3 0.0217
Lser 2 4 0.0000000313
C1 3 4 0.0082
Rpar 3 4 12195.1219512195
.ends 860020380028_8.2mF
*******
.subckt 860020381029_10mF 1 2
Rser 1 3 0.028
Lser 2 4 0.000000025
C1 3 4 0.01
Rpar 3 4 10000
.ends 860020381029_10mF
*******
.subckt 860020381030_12mF 1 2
Rser 1 3 0.022
Lser 2 4 0.000000032
C1 3 4 0.012
Rpar 3 4 8333.33333333333
.ends 860020381030_12mF
*******
.subckt 860020472001_4.7uF 1 2
Rser 1 3 2.2120140088
Lser 2 4 3.130984237E-09
C1 3 4 0.0000047
Rpar 3 4 8333333.33333333
.ends 860020472001_4.7uF
*******
.subckt 860020472002_6.8uF 1 2
Rser 1 3 1.7812436345
Lser 2 4 3.665749892E-09
C1 3 4 0.0000068
Rpar 3 4 8333333.33333333
.ends 860020472002_6.8uF
*******
.subckt 860020472003_10uF 1 2
Rser 1 3 2.09781964725
Lser 2 4 3.11315016E-09
C1 3 4 0.00001
Rpar 3 4 8333333.33333333
.ends 860020472003_10uF
*******
.subckt 860020472004_22uF 1 2
Rser 1 3 0.877349121871
Lser 2 4 4.075442206E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860020472004_22uF
*******
.subckt 860020472005_33uF 1 2
Rser 1 3 0.776103109057
Lser 2 4 4.214627183E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860020472005_33uF
*******
.subckt 860020472006_47uF 1 2
Rser 1 3 0.847012153278
Lser 2 4 4.174130858E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860020472006_47uF
*******
.subckt 860020473007_68uF 1 2
Rser 1 3 0.43
Lser 2 4 0.0000000075
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860020473007_68uF
*******
.subckt 860020473008_100uF 1 2
Rser 1 3 0.445
Lser 2 4 0.00000002
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860020473008_100uF
*******
.subckt 860020473009_120uF 1 2
Rser 1 3 0.46
Lser 2 4 0.00000001962
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860020473009_120uF
*******
.subckt 860020473010_150uF 1 2
Rser 1 3 0.25
Lser 2 4 0.0000000206
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860020473010_150uF
*******
.subckt 860020474011_180uF 1 2
Rser 1 3 0.185
Lser 2 4 0.0000000221
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860020474011_180uF
*******
.subckt 860020474012_220uF 1 2
Rser 1 3 0.2
Lser 2 4 0.0000000202
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860020474012_220uF
*******
.subckt 860020474013_330uF 1 2
Rser 1 3 0.195
Lser 2 4 0.0000000235
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860020474013_330uF
*******
.subckt 860020474014_470uF 1 2
Rser 1 3 0.108
Lser 2 4 0.0000000216
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860020474014_470uF
*******
.subckt 860020475015_560uF 1 2
Rser 1 3 0.133
Lser 2 4 0.0000000272
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860020475015_560uF
*******
.subckt 860020475016_680uF 1 2
Rser 1 3 0.087
Lser 2 4 0.0000000276
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860020475016_680uF
*******
.subckt 860020475017_820uF 1 2
Rser 1 3 0.105
Lser 2 4 0.0000000268
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860020475017_820uF
*******
.subckt 860020475018_1mF 1 2
Rser 1 3 0.086
Lser 2 4 0.0000000268
C1 3 4 0.001
Rpar 3 4 100000
.ends 860020475018_1mF
*******
.subckt 860020478019_1.2mF 1 2
Rser 1 3 0.065
Lser 2 4 0.000000027
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860020478019_1.2mF
*******
.subckt 860020478020_1.5mF 1 2
Rser 1 3 0.0525
Lser 2 4 0.0000000275
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860020478020_1.5mF
*******
.subckt 860020478021_1.8mF 1 2
Rser 1 3 0.044
Lser 2 4 0.000000032
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860020478021_1.8mF
*******
.subckt 860020478022_2.2mF 1 2
Rser 1 3 0.044
Lser 2 4 1.3615768879E-08
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860020478022_2.2mF
*******
.subckt 860020480023_2.7mF 1 2
Rser 1 3 0.043
Lser 2 4 0.0000000341
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860020480023_2.7mF
*******
.subckt 860020480024_3.3mF 1 2
Rser 1 3 0.04
Lser 2 4 0.0000000286
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860020480024_3.3mF
*******
.subckt 860020480025_3.9mF 1 2
Rser 1 3 0.035
Lser 2 4 0.0000000294
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860020480025_3.9mF
*******
.subckt 860020480026_4.7mF 1 2
Rser 1 3 0.03329
Lser 2 4 1.9406012029E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860020480026_4.7mF
*******
.subckt 860020480027_5.6mF 1 2
Rser 1 3 0.0285
Lser 2 4 0.0000000267
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860020480027_5.6mF
*******
.subckt 860020481028_6.8mF 1 2
Rser 1 3 0.029
Lser 2 4 0.000000026
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860020481028_6.8mF
*******
.subckt 860020481029_8.2mF 1 2
Rser 1 3 0.026
Lser 2 4 0.000000032
C1 3 4 0.0082
Rpar 3 4 12195.1219512195
.ends 860020481029_8.2mF
*******
.subckt 860020572001_4.7uF 1 2
Rser 1 3 1.87175337986
Lser 2 4 3.109314535E-09
C1 3 4 0.0000047
Rpar 3 4 11666666.6666667
.ends 860020572001_4.7uF
*******
.subckt 860020572002_6.8uF 1 2
Rser 1 3 2.05012585203
Lser 2 4 2.747361472E-09
C1 3 4 0.0000068
Rpar 3 4 11666666.6666667
.ends 860020572002_6.8uF
*******
.subckt 860020572003_10uF 1 2
Rser 1 3 2.05181792146
Lser 2 4 3.250120717E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860020572003_10uF
*******
.subckt 860020572004_22uF 1 2
Rser 1 3 1.02865081029
Lser 2 4 3.959469941E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 860020572004_22uF
*******
.subckt 860020572005_33uF 1 2
Rser 1 3 0.455999795768
Lser 2 4 4.466402969E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860020572005_33uF
*******
.subckt 860020572006_47uF 1 2
Rser 1 3 0.411275007416
Lser 2 4 4.275625994E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860020572006_47uF
*******
.subckt 860020573007_68uF 1 2
Rser 1 3 0.472327211005
Lser 2 4 4.943461204E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860020573007_68uF
*******
.subckt 860020573008_100uF 1 2
Rser 1 3 0.315
Lser 2 4 0.0000000195
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860020573008_100uF
*******
.subckt 860020574009_120uF 1 2
Rser 1 3 0.407676240681
Lser 2 4 5.414772923E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860020574009_120uF
*******
.subckt 860020574010_150uF 1 2
Rser 1 3 0.187
Lser 2 4 0.0000000259
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860020574010_150uF
*******
.subckt 860020574011_180uF 1 2
Rser 1 3 0.18
Lser 2 4 0.0000000185
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860020574011_180uF
*******
.subckt 860020574012_220uF 1 2
Rser 1 3 0.185
Lser 2 4 0.00000001925
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860020574012_220uF
*******
.subckt 860020575013_330uF 1 2
Rser 1 3 0.135
Lser 2 4 0.000000027
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860020575013_330uF
*******
.subckt 860020575014_470uF 1 2
Rser 1 3 0.098
Lser 2 4 0.0000000208
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860020575014_470uF
*******
.subckt 860020575015_560uF 1 2
Rser 1 3 0.109
Lser 2 4 0.0000000267
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860020575015_560uF
*******
.subckt 860020575016_680uF 1 2
Rser 1 3 0.075
Lser 2 4 0.0000000215
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860020575016_680uF
*******
.subckt 860020578017_820uF 1 2
Rser 1 3 0.066
Lser 2 4 0.0000000283
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860020578017_820uF
*******
.subckt 860020578018_1mF 1 2
Rser 1 3 0.067
Lser 2 4 0.000000024
C1 3 4 0.001
Rpar 3 4 100000
.ends 860020578018_1mF
*******
.subckt 860020578019_1.2mF 1 2
Rser 1 3 0.07
Lser 2 4 0.0000000273
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860020578019_1.2mF
*******
.subckt 860020578020_1.5mF 1 2
Rser 1 3 0.058
Lser 2 4 0.0000000195
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860020578020_1.5mF
*******
.subckt 860020580021_1.8mF 1 2
Rser 1 3 0.045
Lser 2 4 0.0000000301
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860020580021_1.8mF
*******
.subckt 860020580022_2.2mF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000276
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860020580022_2.2mF
*******
.subckt 860020580023_2.7mF 1 2
Rser 1 3 0.0365
Lser 2 4 0.0000000296
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860020580023_2.7mF
*******
.subckt 860020580024_3.3mF 1 2
Rser 1 3 0.028
Lser 2 4 0.000000029
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860020580024_3.3mF
*******
.subckt 860020581025_3.9mF 1 2
Rser 1 3 0.034
Lser 2 4 0.0000000342
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860020581025_3.9mF
*******
.subckt 860020581026_4.7mF 1 2
Rser 1 3 0.03446
Lser 2 4 2.0572094731E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860020581026_4.7mF
*******
.subckt 860020581027_5.6mF 1 2
Rser 1 3 0.027
Lser 2 4 0.0000000361
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860020581027_5.6mF
*******
.subckt 860020672001_100nF 1 2
Rser 1 3 3.11019656901
Lser 2 4 3.825980172E-09
C1 3 4 0.0000001
Rpar 3 4 16666666.6666667
.ends 860020672001_100nF
*******
.subckt 860020672002_220nF 1 2
Rser 1 3 2.48309672257
Lser 2 4 3.190305669E-09
C1 3 4 0.00000022
Rpar 3 4 16666666.6666667
.ends 860020672002_220nF
*******
.subckt 860020672003_330nF 1 2
Rser 1 3 1.81202042505
Lser 2 4 3.525636074E-09
C1 3 4 0.00000033
Rpar 3 4 16666666.6666667
.ends 860020672003_330nF
*******
.subckt 860020672004_470nF 1 2
Rser 1 3 2.68264389854
Lser 2 4 3.497025752E-09
C1 3 4 0.00000047
Rpar 3 4 16666666.6666667
.ends 860020672004_470nF
*******
.subckt 860020672005_1uF 1 2
Rser 1 3 2.33634667339
Lser 2 4 3.377360078E-09
C1 3 4 0.000001
Rpar 3 4 16666666.6666667
.ends 860020672005_1uF
*******
.subckt 860020672006_2.2uF 1 2
Rser 1 3 2.32277177427
Lser 2 4 5.676908907E-09
C1 3 4 0.0000022
Rpar 3 4 16666666.6666667
.ends 860020672006_2.2uF
*******
.subckt 860020672007_3.3uF 1 2
Rser 1 3 1.7619273272
Lser 2 4 3.377157672E-09
C1 3 4 0.0000033
Rpar 3 4 16666666.6666667
.ends 860020672007_3.3uF
*******
.subckt 860020672008_4.7uF 1 2
Rser 1 3 1.81832614741
Lser 2 4 3.00314651E-09
C1 3 4 0.0000047
Rpar 3 4 16666666.6666667
.ends 860020672008_4.7uF
*******
.subckt 860020672009_6.8uF 1 2
Rser 1 3 0.98
Lser 2 4 0.0000000065
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 860020672009_6.8uF
*******
.subckt 860020672010_10uF 1 2
Rser 1 3 1.8698485068
Lser 2 4 3.491870716E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860020672010_10uF
*******
.subckt 860020672011_22uF 1 2
Rser 1 3 0.725557254649
Lser 2 4 4.139560626E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860020672011_22uF
*******
.subckt 860020672012_33uF 1 2
Rser 1 3 0.776398688815
Lser 2 4 3.803472676E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860020672012_33uF
*******
.subckt 860020673013_47uF 1 2
Rser 1 3 0.379063116335
Lser 2 4 5.814672698E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860020673013_47uF
*******
.subckt 860020673014_68uF 1 2
Rser 1 3 0.564800816615
Lser 2 4 4.23651978E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860020673014_68uF
*******
.subckt 860020674015_100uF 1 2
Rser 1 3 0.23
Lser 2 4 0.000000022
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860020674015_100uF
*******
.subckt 860020674016_120uF 1 2
Rser 1 3 0.2
Lser 2 4 0.0000000226
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860020674016_120uF
*******
.subckt 860020675017_120uF 1 2
Rser 1 3 0.215
Lser 2 4 0.0000000227
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860020675017_120uF
*******
.subckt 860020675018_150uF 1 2
Rser 1 3 0.195
Lser 2 4 0.0000000256
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860020675018_150uF
*******
.subckt 860020675019_180uF 1 2
Rser 1 3 0.155
Lser 2 4 0.0000000243
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860020675019_180uF
*******
.subckt 860020675020_220uF 1 2
Rser 1 3 0.195
Lser 2 4 0.0000000194
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860020675020_220uF
*******
.subckt 860020675021_330uF 1 2
Rser 1 3 0.153
Lser 2 4 0.000000018
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860020675021_330uF
*******
.subckt 860020675022_470uF 1 2
Rser 1 3 0.13
Lser 2 4 0.0000000315
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860020675022_470uF
*******
.subckt 860020678023_560uF 1 2
Rser 1 3 0.057
Lser 2 4 0.0000000211
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860020678023_560uF
*******
.subckt 860020678024_680uF 1 2
Rser 1 3 0.055
Lser 2 4 0.0000000215
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860020678024_680uF
*******
.subckt 860020678025_820uF 1 2
Rser 1 3 0.052
Lser 2 4 0.0000000339
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860020678025_820uF
*******
.subckt 860020678026_1mF 1 2
Rser 1 3 0.068
Lser 2 4 0.000000025
C1 3 4 0.001
Rpar 3 4 100000
.ends 860020678026_1mF
*******
.subckt 860020680027_1.2mF 1 2
Rser 1 3 0.038
Lser 2 4 0.0000000302
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860020680027_1.2mF
*******
.subckt 860020680028_1.5mF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000338
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860020680028_1.5mF
*******
.subckt 860020680029_1.8mF 1 2
Rser 1 3 0.03
Lser 2 4 0.0000000325
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860020680029_1.8mF
*******
.subckt 860020680030_2.2mF 1 2
Rser 1 3 0.0295
Lser 2 4 0.0000000301
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860020680030_2.2mF
*******
.subckt 860020681031_2.7mF 1 2
Rser 1 3 0.026
Lser 2 4 0.000000033
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860020681031_2.7mF
*******
.subckt 860020681032_3.3mF 1 2
Rser 1 3 0.031
Lser 2 4 0.0000000285
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860020681032_3.3mF
*******
.subckt 860020772001_100nF 1 2
Rser 1 3 3.13610044602
Lser 2 4 3.808795893E-09
C1 3 4 0.0000001
Rpar 3 4 21000000
.ends 860020772001_100nF
*******
.subckt 860020772002_220nF 1 2
Rser 1 3 2.53725914608
Lser 2 4 3.026158717E-09
C1 3 4 0.00000022
Rpar 3 4 21000000
.ends 860020772002_220nF
*******
.subckt 860020772003_330nF 1 2
Rser 1 3 1.79206812181
Lser 2 4 3.422719259E-09
C1 3 4 0.00000033
Rpar 3 4 21000000
.ends 860020772003_330nF
*******
.subckt 860020772004_470nF 1 2
Rser 1 3 2.4661066526
Lser 2 4 2.836436239E-09
C1 3 4 0.00000047
Rpar 3 4 21000000
.ends 860020772004_470nF
*******
.subckt 860020772005_1uF 1 2
Rser 1 3 2.308284154
Lser 2 4 3.353827633E-09
C1 3 4 0.000001
Rpar 3 4 21000000
.ends 860020772005_1uF
*******
.subckt 860020772006_2.2uF 1 2
Rser 1 3 2.12237009876
Lser 2 4 3.753119462E-09
C1 3 4 0.0000022
Rpar 3 4 21000000
.ends 860020772006_2.2uF
*******
.subckt 860020772007_3.3uF 1 2
Rser 1 3 2.34365396911
Lser 2 4 3.384659869E-09
C1 3 4 0.0000033
Rpar 3 4 21000000
.ends 860020772007_3.3uF
*******
.subckt 860020772008_4.7uF 1 2
Rser 1 3 1.46784557971
Lser 2 4 3.341732332E-09
C1 3 4 0.0000047
Rpar 3 4 21000000
.ends 860020772008_4.7uF
*******
.subckt 860020772009_6.8uF 1 2
Rser 1 3 2.39026815133
Lser 2 4 3.363633194E-09
C1 3 4 0.0000068
Rpar 3 4 14719626.1682243
.ends 860020772009_6.8uF
*******
.subckt 860020772010_10uF 1 2
Rser 1 3 1.67463935163
Lser 2 4 3.765942503E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860020772010_10uF
*******
.subckt 860020773011_22uF 1 2
Rser 1 3 0.413276631743
Lser 2 4 7.120410493E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860020773011_22uF
*******
.subckt 860020773012_33uF 1 2
Rser 1 3 0.71598714939
Lser 2 4 3.513148601E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860020773012_33uF
*******
.subckt 860020773013_47uF 1 2
Rser 1 3 0.464290068005
Lser 2 4 3.776659938E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860020773013_47uF
*******
.subckt 860020774014_68uF 1 2
Rser 1 3 0.175
Lser 2 4 0.0000000087
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860020774014_68uF
*******
.subckt 860020775015_100uF 1 2
Rser 1 3 0.405
Lser 2 4 0.0000000194
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860020775015_100uF
*******
.subckt 860020775016_120uF 1 2
Rser 1 3 0.215
Lser 2 4 0.0000000216
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860020775016_120uF
*******
.subckt 860020775017_150uF 1 2
Rser 1 3 0.129
Lser 2 4 0.0000000243
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860020775017_150uF
*******
.subckt 860020775018_180uF 1 2
Rser 1 3 0.114
Lser 2 4 0.0000000263
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860020775018_180uF
*******
.subckt 860020775019_220uF 1 2
Rser 1 3 0.11
Lser 2 4 0.0000000241
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860020775019_220uF
*******
.subckt 860020778020_330uF 1 2
Rser 1 3 0.071
Lser 2 4 0.0000000265
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860020778020_330uF
*******
.subckt 860020778021_470uF 1 2
Rser 1 3 0.059
Lser 2 4 0.0000000208
C1 3 4 0.00047
Rpar 3 4 212765.957446808
.ends 860020778021_470uF
*******
.subckt 860020778022_560uF 1 2
Rser 1 3 0.09
Lser 2 4 0.0000000318
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860020778022_560uF
*******
.subckt 860020780023_680uF 1 2
Rser 1 3 0.0696
Lser 2 4 0.0000000294
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860020780023_680uF
*******
.subckt 860020780024_820uF 1 2
Rser 1 3 0.059
Lser 2 4 0.000000024
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860020780024_820uF
*******
.subckt 860020780025_1mF 1 2
Rser 1 3 0.027
Lser 2 4 0.0000000267
C1 3 4 0.001
Rpar 3 4 100000
.ends 860020780025_1mF
*******
.subckt 860020780026_1.2mF 1 2
Rser 1 3 0.0305
Lser 2 4 0.0000000333
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860020780026_1.2mF
*******
.subckt 860020781027_1.5mF 1 2
Rser 1 3 0.032
Lser 2 4 0.000000027
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860020781027_1.5mF
*******
.subckt 860021373001_470nF 1 2
Rser 1 3 1.9
Lser 2 4 0.00000000002
C1 3 4 0.00000047
Rpar 3 4 133333333.333333
.ends 860021373001_470nF
*******
.subckt 860021373002_1uF 1 2
Rser 1 3 1.43619741628
Lser 2 4 3.80946011E-09
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 860021373002_1uF
*******
.subckt 860021373003_2.2uF 1 2
Rser 1 3 1.2304311994
Lser 2 4 3.775737786E-09
C1 3 4 0.0000022
Rpar 3 4 45454545.4545455
.ends 860021373003_2.2uF
*******
.subckt 860021373005_3.3uF 1 2
Rser 1 3 1.3222450716
Lser 2 4 5.007147053E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 860021373005_3.3uF
*******
.subckt 860021373025_4.7uF 1 2
Rser 1 3 0.84
Lser 2 4 0.000000000019
C1 3 4 0.0000047
Rpar 3 4 7092198.58156028
.ends 860021373025_4.7uF
*******
.subckt 860021374004_2.2uF 1 2
Rser 1 3 1.40205839386
Lser 2 4 4.772007064E-09
C1 3 4 0.0000022
Rpar 3 4 45454545.4545455
.ends 860021374004_2.2uF
*******
.subckt 860021374006_3.3uF 1 2
Rser 1 3 0.989809251237
Lser 2 4 4.107108381E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 860021374006_3.3uF
*******
.subckt 860021374008_4.7uF 1 2
Rser 1 3 0.780247662714
Lser 2 4 3.621111012E-09
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 860021374008_4.7uF
*******
.subckt 860021374009_6.8uF 1 2
Rser 1 3 0.830156310587
Lser 2 4 5.0462049E-09
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 860021374009_6.8uF
*******
.subckt 860021375007_3.3uF 1 2
Rser 1 3 1.25878201217
Lser 2 4 4.014372865E-09
C1 3 4 0.0000033
Rpar 3 4 30303030.3030303
.ends 860021375007_3.3uF
*******
.subckt 860021375010_6.8uF 1 2
Rser 1 3 0.733913311919
Lser 2 4 4.417511372E-09
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 860021375010_6.8uF
*******
.subckt 860021375011_10uF 1 2
Rser 1 3 0.611701901159
Lser 2 4 4.242583346E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860021375011_10uF
*******
.subckt 860021375012_22uF 1 2
Rser 1 3 0.408321609223
Lser 2 4 4.41071527E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860021375012_22uF
*******
.subckt 860021378013_22uF 1 2
Rser 1 3 0.595071057581
Lser 2 4 6.825738473E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860021378013_22uF
*******
.subckt 860021378014_33uF 1 2
Rser 1 3 0.411039493813
Lser 2 4 6.048850153E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860021378014_33uF
*******
.subckt 860021380015_47uF 1 2
Rser 1 3 0.60266
Lser 2 4 1.4438885117E-08
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860021380015_47uF
*******
.subckt 860021380016_56uF 1 2
Rser 1 3 0.480680508203
Lser 2 4 1.2229475031E-08
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860021380016_56uF
*******
.subckt 860021380017_68uF 1 2
Rser 1 3 0.475658642144
Lser 2 4 1.3386184191E-08
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860021380017_68uF
*******
.subckt 860021380018_82uF 1 2
Rser 1 3 0.404141160298
Lser 2 4 1.1207183067E-08
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860021380018_82uF
*******
.subckt 860021380020_100uF 1 2
Rser 1 3 0.358015810583
Lser 2 4 1.0964407714E-08
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860021380020_100uF
*******
.subckt 860021381019_82uF 1 2
Rser 1 3 0.440713489779
Lser 2 4 1.2672547142E-08
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860021381019_82uF
*******
.subckt 860021381021_120uF 1 2
Rser 1 3 0.365395489766
Lser 2 4 1.2562615098E-08
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860021381021_120uF
*******
.subckt 860021381022_150uF 1 2
Rser 1 3 0.292087676123
Lser 2 4 1.0796501344E-08
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860021381022_150uF
*******
.subckt 860021381024_180uF 1 2
Rser 1 3 0.255822762362
Lser 2 4 9.144474952E-09
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860021381024_180uF
*******
.subckt 860021383023_150uF 1 2
Rser 1 3 0.312793214947
Lser 2 4 1.1479296572E-08
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860021383023_150uF
*******
.subckt 860020684033_10mF 1 2
Rser 1 3 0.0177
Lser 2 4 0.0000000226
C1 3 4 0.01
Rpar 3 4 10000
.ends 860020684033_10mF
*******
.subckt 860021374027_22uF 1 2
Rser 1 3 0.44
Lser 2 4 0.00000000001
C1 3 4 0.000022
Rpar 3 4 1515151.51515152
.ends 860021374027_22uF
*******
