**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-AT1H
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 860240272001_47uF 1 2
Rser 1 3 1.40169642531
Lser 2 4 3.871861968E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860240272001_47uF
*******
.subckt 860240272002_68uF 1 2
Rser 1 3 1.45957602277
Lser 2 4 5.564041279E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860240272002_68uF
*******
.subckt 860240273003_100uF 1 2
Rser 1 3 0.55
Lser 2 4 0.0000000035
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860240273003_100uF
*******
.subckt 860240273004_150uF 1 2
Rser 1 3 0.47
Lser 2 4 4.622534653E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860240273004_150uF
*******
.subckt 860240273005_220uF 1 2
Rser 1 3 0.5
Lser 2 4 4.103221197E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860240273005_220uF
*******
.subckt 860240274006_330uF 1 2
Rser 1 3 0.25
Lser 2 4 0.0000000012
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860240274006_330uF
*******
.subckt 860240275007_470uF 1 2
Rser 1 3 0.19
Lser 2 4 0.0000000015
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860240275007_470uF
*******
.subckt 860240275008_1mF 1 2
Rser 1 3 0.093
Lser 2 4 0.0000000019
C1 3 4 0.001
Rpar 3 4 100000
.ends 860240275008_1mF
*******
.subckt 860240278009_2.2mF 1 2
Rser 1 3 0.057
Lser 2 4 0.0000000035
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860240278009_2.2mF
*******
.subckt 860240280010_3.3mF 1 2
Rser 1 3 0.043
Lser 2 4 4.76579264672459E-09
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860240280010_3.3mF
*******
.subckt 860240372001_33uF 1 2
Rser 1 3 1.45287605459
Lser 2 4 3.252512554E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860240372001_33uF
*******
.subckt 860240372002_47uF 1 2
Rser 1 3 1.23739536051
Lser 2 4 3.513901242E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860240372002_47uF
*******
.subckt 860240373003_68uF 1 2
Rser 1 3 0.910878310644
Lser 2 4 4.03203322E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860240373003_68uF
*******
.subckt 860240374004_100uF 1 2
Rser 1 3 0.346593548429
Lser 2 4 4.16242534E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860240374004_100uF
*******
.subckt 860240374005_150uF 1 2
Rser 1 3 0.477911623357
Lser 2 4 4.128536017E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860240374005_150uF
*******
.subckt 860240374006_220uF 1 2
Rser 1 3 0.232
Lser 2 4 0.0000000015
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860240374006_220uF
*******
.subckt 860240374007_330uF 1 2
Rser 1 3 0.175
Lser 2 4 0.0000000025
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860240374007_330uF
*******
.subckt 860240375008_470uF 1 2
Rser 1 3 0.137
Lser 2 4 0.000000002
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860240375008_470uF
*******
.subckt 860240378009_1mF 1 2
Rser 1 3 0.071
Lser 2 4 0.0000000055
C1 3 4 0.001
Rpar 3 4 100000
.ends 860240378009_1mF
*******
.subckt 860240380010_2.2mF 1 2
Rser 1 3 0.039
Lser 2 4 0.0000000075
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860240380010_2.2mF
*******
.subckt 860240472001_22uF 1 2
Rser 1 3 1.41461577405
Lser 2 4 5.415005782E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860240472001_22uF
*******
.subckt 860240472002_33uF 1 2
Rser 1 3 1.26000876057
Lser 2 4 3.636367687E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860240472002_33uF
*******
.subckt 860240473003_47uF 1 2
Rser 1 3 0.716766005667
Lser 2 4 4.300549436E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860240473003_47uF
*******
.subckt 860240474004_68uF 1 2
Rser 1 3 0.359211639719
Lser 2 4 4.499207576E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860240474004_68uF
*******
.subckt 860240474005_100uF 1 2
Rser 1 3 0.315
Lser 2 4 0.0000000013
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860240474005_100uF
*******
.subckt 860240475006_150uF 1 2
Rser 1 3 0.172
Lser 2 4 0.000000003
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860240475006_150uF
*******
.subckt 860240475007_220uF 1 2
Rser 1 3 0.27
Lser 2 4 0.0000000221
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860240475007_220uF
*******
.subckt 860240475008_330uF 1 2
Rser 1 3 0.112
Lser 2 4 0.0000000035
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860240475008_330uF
*******
.subckt 860240475009_470uF 1 2
Rser 1 3 0.09
Lser 2 4 0.000000005
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860240475009_470uF
*******
.subckt 860240478010_1mF 1 2
Rser 1 3 0.05
Lser 2 4 0.00000001
C1 3 4 0.001
Rpar 3 4 100000
.ends 860240478010_1mF
*******
.subckt 860240480011_2.2mF 1 2
Rser 1 3 0.036
Lser 2 4 0.0000000055
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860240480011_2.2mF
*******
.subckt 860240572001_10uF 1 2
Rser 1 3 0.9
Lser 2 4 3.044427204E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860240572001_10uF
*******
.subckt 860240572002_22uF 1 2
Rser 1 3 1.33849819282
Lser 2 4 3.216545731E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 860240572002_22uF
*******
.subckt 860240573003_33uF 1 2
Rser 1 3 0.783576881536
Lser 2 4 4.861643715E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860240573003_33uF
*******
.subckt 860240574004_47uF 1 2
Rser 1 3 0.682883081334
Lser 2 4 4.912250742E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860240574004_47uF
*******
.subckt 860240574005_68uF 1 2
Rser 1 3 0.3907341567
Lser 2 4 5.089062183E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860240574005_68uF
*******
.subckt 860240575006_100uF 1 2
Rser 1 3 0.235
Lser 2 4 0.000000003
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860240575006_100uF
*******
.subckt 860240575007_150uF 1 2
Rser 1 3 0.18
Lser 2 4 0.000000003
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860240575007_150uF
*******
.subckt 860240575008_220uF 1 2
Rser 1 3 0.125
Lser 2 4 0.0000000045
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860240575008_220uF
*******
.subckt 860240578009_330uF 1 2
Rser 1 3 0.092
Lser 2 4 0.000000007
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860240578009_330uF
*******
.subckt 860240578010_470uF 1 2
Rser 1 3 0.082
Lser 2 4 0.000000007
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860240578010_470uF
*******
.subckt 860240580011_1mF 1 2
Rser 1 3 0.041
Lser 2 4 0.000000009
C1 3 4 0.001
Rpar 3 4 100000
.ends 860240580011_1mF
*******
.subckt 860240672001_6.8uF 1 2
Rser 1 3 1.369893426
Lser 2 4 3.660038331E-09
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 860240672001_6.8uF
*******
.subckt 860240672002_10uF 1 2
Rser 1 3 1.96224521591
Lser 2 4 4.356061895E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860240672002_10uF
*******
.subckt 860240673003_22uF 1 2
Rser 1 3 0.721604412351
Lser 2 4 3.657813236E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860240673003_22uF
*******
.subckt 860240674004_33uF 1 2
Rser 1 3 0.24
Lser 2 4 0.000000005
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860240674004_33uF
*******
.subckt 860240674005_47uF 1 2
Rser 1 3 0.38172487193
Lser 2 4 4.210500451E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860240674005_47uF
*******
.subckt 860240675006_68uF 1 2
Rser 1 3 0.272
Lser 2 4 0.0000000032
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860240675006_68uF
*******
.subckt 860240675007_100uF 1 2
Rser 1 3 0.22306
Lser 2 4 9.472671859E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860240675007_100uF
*******
.subckt 860240675008_150uF 1 2
Rser 1 3 0.141
Lser 2 4 0.000000006
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860240675008_150uF
*******
.subckt 860240678009_220uF 1 2
Rser 1 3 0.12295
Lser 2 4 1.1548923515E-08
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860240678009_220uF
*******
.subckt 860240678010_330uF 1 2
Rser 1 3 0.079
Lser 2 4 9.15240353855245E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860240678010_330uF
*******
.subckt 860240680011_470uF 1 2
Rser 1 3 0.048
Lser 2 4 0.000000009
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860240680011_470uF
*******
.subckt 860240681012_1mF 1 2
Rser 1 3 0.036
Lser 2 4 0.00000001
C1 3 4 0.001
Rpar 3 4 100000
.ends 860240681012_1mF
*******
.subckt 860240975001_10uF 1 2
Rser 1 3 0.6
Lser 2 4 0.33934242
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860240975001_10uF
*******
.subckt 860240975002_22uF 1 2
Rser 1 3 0.719871933466
Lser 2 4 4.565216798E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 860240975002_22uF
*******
.subckt 860240978003_33uF 1 2
Rser 1 3 0.3
Lser 2 4 4.884412961E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860240978003_33uF
*******
.subckt 860240978004_47uF 1 2
Rser 1 3 0.448655216894
Lser 2 4 6.431602964E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860240978004_47uF
*******
.subckt 860240978005_68uF 1 2
Rser 1 3 0.324160550936
Lser 2 4 6.58149596E-09
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860240978005_68uF
*******
.subckt 860240981006_100uF 1 2
Rser 1 3 0.241099978468
Lser 2 4 1.0399106109E-08
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860240981006_100uF
*******
.subckt 860240981007_150uF 1 2
Rser 1 3 0.13
Lser 2 4 1.1041262827E-08
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860240981007_150uF
*******
.subckt 860240981008_220uF 1 2
Rser 1 3 0.146888860269
Lser 2 4 1.4561098727E-08
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860240981008_220uF
*******
.subckt 860241075003_10uF 1 2
Rser 1 3 0.73654396039
Lser 2 4 4.498665017E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860241075003_10uF
*******
.subckt 860241075004_22uF 1 2
Rser 1 3 0.619580383999
Lser 2 4 4.370805351E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860241075004_22uF
*******
.subckt 860241078002_47uF 1 2
Rser 1 3 0.34485838389
Lser 2 4 4.950182861E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860241078002_47uF
*******
.subckt 860241078005_33uF 1 2
Rser 1 3 0.506188561351
Lser 2 4 7.156208262E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860241078005_33uF
*******
.subckt 860241080006_68uF 1 2
Rser 1 3 0.261171828785
Lser 2 4 0.000000013546
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860241080006_68uF
*******
.subckt 860241081001_330uF 1 2
Rser 1 3 0.129477441882
Lser 2 4 1.0036580705E-08
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860241081001_330uF
*******
.subckt 860241081007_100uF 1 2
Rser 1 3 0.18
Lser 2 4 8.821406195E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860241081007_100uF
*******
.subckt 860241081008_150uF 1 2
Rser 1 3 0.16839264055
Lser 2 4 1.3355271602E-08
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860241081008_150uF
*******
.subckt 860241081009_220uF 1 2
Rser 1 3 0.113285691859
Lser 2 4 1.1535560401E-08
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860241081009_220uF
*******
.subckt 860241175001_10uF 1 2
Rser 1 3 0.7
Lser 2 4 0.00000001
C1 3 4 0.00001
Rpar 3 4 1600000
.ends 860241175001_10uF
*******
.subckt 860241175002_22uF 1 2
Rser 1 3 0.3
Lser 2 4 4.908482481E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860241175002_22uF
*******
.subckt 860241178002_22uF 1 2
Rser 1 3 1.6
Lser 2 4 0.000000007
C1 3 4 0.000022
Rpar 3 4 1531250
.ends 860241178002_22uF
*******
.subckt 860241178003_33uF 1 2
Rser 1 3 1.2
Lser 2 4 0.000000006495
C1 3 4 0.000033
Rpar 3 4 1744186.04651163
.ends 860241178003_33uF
*******
.subckt 860241180004_47uF 1 2
Rser 1 3 0.276875722098
Lser 2 4 1.0521240941E-08
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860241180004_47uF
*******
.subckt 860241181005_68uF 1 2
Rser 1 3 0.225510181399
Lser 2 4 1.2339052472E-08
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860241181005_68uF
*******
.subckt 860241181006_100uF 1 2
Rser 1 3 0.208676890185
Lser 2 4 1.4288872982E-08
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860241181006_100uF
*******
.subckt 860241181007_150uF 1 2
Rser 1 3 0.223518441256
Lser 2 4 1.1835999533E-08
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860241181007_150uF
*******
.subckt 860241375001_6.8uF 1 2
Rser 1 3 0.743001817068
Lser 2 4 4.687155572E-09
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 860241375001_6.8uF
*******
.subckt 860241375002_10uF 1 2
Rser 1 3 0.652367911032
Lser 2 4 4.404273931E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860241375002_10uF
*******
.subckt 860241378003_22uF 1 2
Rser 1 3 0.5269419234
Lser 2 4 7.545296913E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860241378003_22uF
*******
.subckt 860241380015_47uF 1 2
Rser 1 3 0.3
Lser 2 4 0.000000008
C1 3 4 0.000047
Rpar 3 4 1408450.70422535
.ends 860241380015_47uF
*******
.subckt 860241381004_33uF 1 2
Rser 1 3 0.592971221632
Lser 2 4 1.047241225E-08
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860241381004_33uF
*******
.subckt 860241381005_47uF 1 2
Rser 1 3 0.52487507871
Lser 2 4 1.2008960083E-08
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860241381005_47uF
*******
.subckt 860241381006_68uF 1 2
Rser 1 3 0.27
Lser 2 4 0.00000001
C1 3 4 0.000068
Rpar 3 4 1228956.22895623
.ends 860241381006_68uF
*******
.subckt 860241381008_82uF 1 2
Rser 1 3 0.25
Lser 2 4 0.000000008
C1 3 4 0.000082
Rpar 3 4 1083569.40509915
.ends 860241381008_82uF
*******
.subckt 860241478002_6.8uF 1 2
Rser 1 3 0.86431
Lser 2 4 9.87132149E-09
C1 3 4 0.0000068
Rpar 3 4 14705882.3529412
.ends 860241478002_6.8uF
*******
.subckt 860241478003_10uF 1 2
Rser 1 3 1.01763676485
Lser 2 4 9.918160074E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860241478003_10uF
*******
.subckt 860241478004_22uF 1 2
Rser 1 3 0.69929
Lser 2 4 1.0635926305E-08
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860241478004_22uF
*******
.subckt 860241480001_100uF 1 2
Rser 1 3 0.37418
Lser 2 4 1.3712726643E-08
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860241480001_100uF
*******
.subckt 860241480005_22uF 1 2
Rser 1 3 0.75671
Lser 2 4 1.3090545796E-08
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860241480005_22uF
*******
.subckt 860241481006_33uF 1 2
Rser 1 3 0.61935
Lser 2 4 1.3714343001E-08
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860241481006_33uF
*******
.subckt 860241481007_47uF 1 2
Rser 1 3 0.54293
Lser 2 4 1.3955585143E-08
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860241481007_47uF
*******
