**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  SMT Full-color Side View Waterclear 
* Matchcode:              WL-SFSW
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Ella      
* Date and Time:          2022-11-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1204_155124M173200 1 2 3 4 
D1 1 2 Blue
.MODEL Blue D
+ IS=24.280E-12
+ N=3.8516
+ RS=1.1745
+ IKF=792.64E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
+ TT=5.0000E-9
D2 1 3 Green
.MODEL Green D
+ IS=118.19E-18
+ N=3.0436
+ RS=.43217
+ IKF=722.66E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
+ TT=5.0000E-9
D3 1 4 Red
.MODEL Red D
+ IS=10.000E-21
+ N=1.7618
+ RS=1.0000E-6
+ IKF=2.0622E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 1204_155124M173200A 1 2 3 4 
D1 4 1 Green
.MODEL Green D
+ IS=847.93E-18
+ N=3.4400
+ RS=.51865
+ IKF=753.31E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
+ TT=5.0000E-9
D2 4 2 Red
.MODEL Red D
+ IS=10.000E-21
+ N=1.7618
+ RS=1.0000E-6
+ IKF=2.0622E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
+ TT=5.0000E-9
D3 4 3 Blue
.MODEL Blue D
+ IS=209.14E-15
+ N=4.2784
+ RS=.78026
+ IKF=865.02E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=1.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 1204_155124M172400 1 2 3 4 
D1 1 2 Blue
.MODEL Blue D
+ IS=1.4711E-15
+ N=3.3923
+ RS=.54588
+ IKF=413.48E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
D2 1 3 Green
.MODEL Green D
+ IS=7.2379E-15
+ N=3.3919
+ RS=.54629
+ IKF=413.19E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
D3 1 4 Red
.MODEL Red D
+ IS=10.010E-21
+ N=1.9114
+ RS=1.0000E-6
+ IKF=47.488E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ TT=5.0000E-9
.ends
******
























