**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  Power Molded Flatwire Inductor
* Matchcode:              WE-PMFI
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          2/12/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 201610_74479320165110_0.1u 1 2
Rp 1 2 283.9412
Cp 1 2 2.412999p
Rs 1 N3 0.0072
L1 N3 2 0.0997761u
.ends 201610_74479320165110_0.1u
*******
.subckt 201610_74479320165124_0.24u 1 2
Rp 1 2 415.4765
Cp 1 2 4.5849p
Rs 1 N3 0.0105
L1 N3 2 0.2331993u
.ends 201610_74479320165124_0.24u
*******
.subckt 201610_74479320165133_0.33u 1 2
Rp 1 2 516.452
Cp 1 2 4.0599p
Rs 1 N3 0.0151
L1 N3 2 0.2980548u
.ends 201610_74479320165133_0.33u
*******
.subckt 201610_74479320165147_0.47u 1 2
Rp 1 2 548.1689
Cp 1 2 5.7371p
Rs 1 N3 0.0184
L1 N3 2 0.4392495u
.ends 201610_74479320165147_0.47u
*******
.subckt 201610_74479320165168_0.68u 1 2
Rp 1 2 840.6128
Cp 1 2 5.0718p
Rs 1 N3 0.0248
L1 N3 2 0.6142667u
.ends 201610_74479320165168_0.68u
*******
.subckt 201610_74479320165210_1u 1 2
Rp 1 2 781.0979
Cp 1 2 6.3458p
Rs 1 N3 0.0317
L1 N3 2 0.9017093u
.ends 201610_74479320165210_1u
*******
.subckt 201610_74479320165215_1.5u 1 2
Rp 1 2 1365
Cp 1 2 5.8292p
Rs 1 N3 0.0561
L1 N3 2 1.4699u
.ends 201610_74479320165215_1.5u
*******
.subckt 201610_74479320165222_2.2u 1 2
Rp 1 2 2347
Cp 1 2 4.8687p
Rs 1 N3 0.0819
L1 N3 2 1.985u
.ends 201610_74479320165222_2.2u
*******
.subckt 201610_74479320165233_3.3u 1 2
Rp 1 2 2754.9
Cp 1 2 6.3111p
Rs 1 N3 0.146
L1 N3 2 3.3817u
.ends 201610_74479320165233_3.3u
*******
.subckt 201610_74479320165247_4.7u 1 2
Rp 1 2 3169.2
Cp 1 2 6.5249p
Rs 1 N3 0.195
L1 N3 2 4.4961u
.ends 201610_74479320165247_4.7u
*******
.subckt 201610_74479320165268_6.8u 1 2
Rp 1 2 5125.71428571429
Cp 1 2 5.3254p
Rs 1 N3 0.458
L1 N3 2 6.242u
.ends 201610_74479320165268_6.8u
*******
.subckt 252012_74479325207110_0.1u 1 2
Rp 1 2 210.569
Cp 1 2 2.0186995p
Rs 1 N3 0.0056
L1 N3 2 0.0659748u
.ends 252012_74479325207110_0.1u
*******
.subckt 252012_74479325207124_0.24u 1 2
Rp 1 2 552.5746
Cp 1 2 4.008p
Rs 1 N3 0.0111
L1 N3 2 0.2302043u
.ends 252012_74479325207124_0.24u
*******
.subckt 252012_74479325207133_0.33u 1 2
Rp 1 2 426.3608
Cp 1 2 5.5322p
Rs 1 N3 0.0105
L1 N3 2 0.3095u
.ends 252012_74479325207133_0.33u
*******
.subckt 252012_74479325207147_0.47u 1 2
Rp 1 2 537.0959
Cp 1 2 5.9841p
Rs 1 N3 0.0113
L1 N3 2 0.4494777u
.ends 252012_74479325207147_0.47u
*******
.subckt 252012_74479325207168_0.68u 1 2
Rp 1 2 678.4212
Cp 1 2 8.2081p
Rs 1 N3 0.0153
L1 N3 2 0.6149067u
.ends 252012_74479325207168_0.68u
*******
.subckt 252012_74479325207210_1u 1 2
Rp 1 2 1030.5355
Cp 1 2 7.7965p
Rs 1 N3 0.0238
L1 N3 2 0.9752471u
.ends 252012_74479325207210_1u
*******
.subckt 252012_74479325207215_1.5u 1 2
Rp 1 2 1669.6
Cp 1 2 8.1081p
Rs 1 N3 0.0373
L1 N3 2 1.5056u
.ends 252012_74479325207215_1.5u
*******
.subckt 252012_74479325207222_2.2u 1 2
Rp 1 2 1982.7
Cp 1 2 7.9778p
Rs 1 N3 0.0501
L1 N3 2 2.0781u
.ends 252012_74479325207222_2.2u
*******
.subckt 252012_74479325207233_3.3u 1 2
Rp 1 2 2667.9
Cp 1 2 9.3574p
Rs 1 N3 0.0848
L1 N3 2 3.0036u
.ends 252012_74479325207233_3.3u
*******
.subckt 252012_74479325207247_4.7u 1 2
Rp 1 2 3182.9
Cp 1 2 9.0759p
Rs 1 N3 0.114
L1 N3 2 4.6455u
.ends 252012_74479325207247_4.7u
*******
.subckt 252012_74479325207268_6.8u 1 2
Rp 1 2 3805.4
Cp 1 2 7.617p
Rs 1 N3 0.205
L1 N3 2 6.1708u
.ends 252012_74479325207268_6.8u
*******
.subckt 322512_74479332257110_0.1u 1 2
Rp 1 2 262.0234
Cp 1 2 1.6953312p
Rs 1 N3 0.0074
L1 N3 2 0.0918745u
.ends 322512_74479332257110_0.1u
*******
.subckt 322512_74479332257124_0.24u 1 2
Rp 1 2 410.4631
Cp 1 2 2.668p
Rs 1 N3 0.0106
L1 N3 2 0.1887002u
.ends 322512_74479332257124_0.24u
*******
.subckt 322512_74479332257133_0.33u 1 2
Rp 1 2 925.5003
Cp 1 2 4.178p
Rs 1 N3 0.0144
L1 N3 2 0.3155138u
.ends 322512_74479332257133_0.33u
*******
.subckt 322512_74479332257147_0.47u 1 2
Rp 1 2 448.4743
Cp 1 2 3.6323p
Rs 1 N3 0.0142
L1 N3 2 0.4449967u
.ends 322512_74479332257147_0.47u
*******
.subckt 322512_74479332257168_0.68u 1 2
Rp 1 2 623.093
Cp 1 2 5.1108p
Rs 1 N3 0.0177
L1 N3 2 0.5806713u
.ends 322512_74479332257168_0.68u
*******
.subckt 322512_74479332257210_1u 1 2
Rp 1 2 908.0213
Cp 1 2 6.5025p
Rs 1 N3 0.0233
L1 N3 2 0.8795647u
.ends 322512_74479332257210_1u
*******
.subckt 322512_74479332257215_1.5u 1 2
Rp 1 2 1229.7
Cp 1 2 6.9957p
Rs 1 N3 0.0365
L1 N3 2 1.38982u
.ends 322512_74479332257215_1.5u
*******
.subckt 322512_74479332257222_2.2u 1 2
Rp 1 2 1612.5
Cp 1 2 6.706p
Rs 1 N3 0.0496
L1 N3 2 1.9717u
.ends 322512_74479332257222_2.2u
*******
.subckt 322512_74479332257233_3.3u 1 2
Rp 1 2 1873.3
Cp 1 2 6.9902p
Rs 1 N3 0.0777
L1 N3 2 3.1365u
.ends 322512_74479332257233_3.3u
*******
.subckt 322512_74479332257247_4.7u 1 2
Rp 1 2 2444.8
Cp 1 2 8.7219p
Rs 1 N3 0.107
L1 N3 2 4.6533u
.ends 322512_74479332257247_4.7u
*******
.subckt 322512_74479332257268_6.8u 1 2
Rp 1 2 4137.8
Cp 1 2 8.5869p
Rs 1 N3 0.17
L1 N3 2 6.5472u
.ends 322512_74479332257268_6.8u
*******
.subckt 353220_74479335329110_0.1u 1 2
Rp 1 2 244.7095
Cp 1 2 2.7559p
Rs 1 N3 0.0048
L1 N3 2 0.0964471u
.ends 353220_74479335329110_0.1u
*******
.subckt 353220_74479335329124_0.24u 1 2
Rp 1 2 402.0035
Cp 1 2 4.6404p
Rs 1 N3 0.0064
L1 N3 2 0.1990607u
.ends 353220_74479335329124_0.24u
*******
.subckt 353220_74479335329133_0.33u 1 2
Rp 1 2 504.9665
Cp 1 2 5.633p
Rs 1 N3 0.0093
L1 N3 2 0.302776u
.ends 353220_74479335329133_0.33u
*******
.subckt 353220_74479335329147_0.47u 1 2
Rp 1 2 712.4074
Cp 1 2 6.2406p
Rs 1 N3 0.0127
L1 N3 2 0.4823098u
.ends 353220_74479335329147_0.47u
*******
.subckt 353220_74479335329168_0.68u 1 2
Rp 1 2 1258.6
Cp 1 2 6.6209p
Rs 1 N3 0.015
L1 N3 2 0.733328u
.ends 353220_74479335329168_0.68u
*******
.subckt 353220_74479335329210_1u 1 2
Rp 1 2 1401.9
Cp 1 2 8.0074p
Rs 1 N3 0.0184
L1 N3 2 1.0162148u
.ends 353220_74479335329210_1u
*******
.subckt 353220_74479335329215_1.5u 1 2
Rp 1 2 1621.1
Cp 1 2 9.42p
Rs 1 N3 0.0253
L1 N3 2 1.6319u
.ends 353220_74479335329215_1.5u
*******
.subckt 353220_74479335329222_2.2u 1 2
Rp 1 2 2535.2
Cp 1 2 10.9292p
Rs 1 N3 0.0316
L1 N3 2 2.3833u
.ends 353220_74479335329222_2.2u
*******
.subckt 353220_74479335329233_3.3u 1 2
Rp 1 2 3922.7
Cp 1 2 10.7255p
Rs 1 N3 0.0529
L1 N3 2 3.6816u
.ends 353220_74479335329233_3.3u
*******
.subckt 353220_74479335329247_4.7u 1 2
Rp 1 2 3860
Cp 1 2 12.4106p
Rs 1 N3 0.0632
L1 N3 2 4.6426u
.ends 353220_74479335329247_4.7u
*******
.subckt 353220_74479335329268_6.8u 1 2
Rp 1 2 4566.5
Cp 1 2 10.4259p
Rs 1 N3 0.118
L1 N3 2 6.9739u
.ends 353220_74479335329268_6.8u
*******
