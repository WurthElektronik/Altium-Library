**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Wirewound Ferrite Bead
* Matchcode:              WE-RFI 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-07-08
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0805A_744760247A_0.47u 1 2
C1 1 N7 159.5136f
L1 1 N1 450n
L2 N1 N2 20.2094n
L3 N2 N3 18.6247n
L4 N3 N4 583.9523p
L5 N4 N5 9.5844n
L6 N5 N6 1.0575
R1 2 N1 6.1204
R2 2 N2 1.0575
R3 2 N3 9.4334
R4 2 N4 287.0525m
R5 2 N5 8.8470
R6 2 N6 7.1327
R7 2 N7 647.9627
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760256A_0.56u 1 2
C1 1 N7 153.5612f
L1 1 N1 530n
L2 N1 N2 26.8088n
L3 N2 N3 20.2434n
L4 N3 N4 584.2412p
L5 N4 N5 9.5854n
L6 N5 N6 2.4030n
R1 2 N1 6.1191
R2 2 N2 1.0634
R3 2 N3 9.4334
R4 2 N4 294.2585m
R5 2 N5 8.8470
R6 2 N6 7.1327
R7 2 N7 647.5479
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760268A_0.68u 1 2
C1 1 N7 136.6774f
L1 1 N1 663.5n
L2 N1 N2 42.4299n
L3 N2 N3 7.5466n
L4 N3 N4 413.2899p
L5 N4 N5 98.1445n
L6 N5 N6 2.5968n
R1 2 N1 9.4018
R2 2 N2 3.2364
R3 2 N3 9.5397
R4 2 N4 3.3780
R5 2 N5 7.2689
R6 2 N6 8.0843
R7 2 N7 841.5979
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760282A_0.82u 1 2
C1 1 N7 138.9514f
L1 1 N1 770n
L2 N1 N2 8.1508n
L3 N2 N3 2.5651n
L4 N3 N4 40.7889n
L5 N4 N5 14.0322n
L6 N5 N6 12.2484n
R1 2 N1 35.1686
R2 2 N2 18.4937
R3 2 N3 21.2775
R4 2 N4 1.3639
R5 2 N5 9.4796
R6 2 N6 8.0236
R7 2 N7 644.7885
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760310A_1u 1 2
C1 1 N7 127.1422f
L1 1 N1 950n
L2 N1 N2 26.8186n
L3 N2 N3 2.9875n
L4 N3 N4 49.6184n
L5 N4 N5 32.3062n
L6 N5 N6 22.7513n
R1 2 N1 35.2122
R2 2 N2 18.5686
R3 2 N3 21.3253
R4 2 N4 2.5096
R5 2 N5 9.4651
R6 2 N6 7.9994
R7 2 N7 642.5452
R8 2 1 10g
.ends
*******
.subckt 0805A_744760312A_1.2u 1 2
C1 1 N7 127.5473f
L1 1 N1 1.15u
L2 N1 N2 33.5362n
L3 N2 N3 2.6037n
L4 N3 N4 41.1788n
L5 N4 N5 61.5148n
L6 N5 N6 29.7561n
R1 2 N1 37.1888
R2 2 N2 17.7304
R3 2 N3 20.6893
R4 2 N4 2.6032
R5 2 N5 9.4682
R6 2 N6 7.9975
R7 2 N7 697.2085
R8 2 1 10g
.ends 
******* 
.subckt 0805A_744760315A_1.5u 1 2
C1 1 N7 123.1843f
L1 1 N1 1.3757u
L2 N1 N2 57.6285n
L3 N2 N3 3.5418n
L4 N3 N4 55.0942n
L5 N4 N5 49.7480n
L6 N5 N6 31.5411n
R1 2 N1 33.7177
R2 2 N2 20.6069
R3 2 N3 22.8943
R4 2 N4 6.4423
R5 2 N5 9.4804
R6 2 N6 8.0146
R7 2 N7 553.8673
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760318A_1.8u 1 2
C1 1 N7 133.8760f
L1 1 N1 1.65u
L2 N1 N2 65.6086n
L3 N2 N3 3.1064n
L4 N3 N4 60.6754n
L5 N4 N5 79.8796n
L6 N5 N6 40.7869n
R1 2 N1 36.1006
R2 2 N2 21.3755
R3 2 N3 23.5436
R4 2 N4 13.1875
R5 2 N5 9.5493
R6 2 N6 8.1022
R7 2 N7 423.1638
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760322A_2.2u 1 2
C1 1 N7 189.8719f
L1 1 N1 1.8u
L2 N1 N2 450.0742n
L3 N2 N3 2.5035n
L4 N3 N4 5.9638n
L5 N4 N5 7.9713n
L6 N5 N6 4.0616n
R1 2 N1 190.9297
R2 2 N2 24.7252
R3 2 N3 25.7638
R4 2 N4 9.0673
R5 2 N5 9.5964
R6 2 N6 8.1937
R7 2 N7 923.0878
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760327A_2.7u 1 2
C1 1 N7 135.9031f
L1 1 N1 2.25u
L2 N1 N2 583.7325n
L3 N2 N3 3.1043n
L4 N3 N4 6.3162n
L5 N4 N5 8.1769n
L6 N5 N6 4.3153n
R1 2 N1 171.6405
R2 2 N2 24.4242
R3 2 N3 25.4783
R4 2 N4 9.0386
R5 2 N5 9.5704
R6 2 N6 8.1571
R7 2 N7 1.4363k
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760333A_3.3u 1 2
C1 1 N7 158.0233f
L1 1 N1 2.8u
L2 N1 N2 619.9642n
L3 N2 N3 750.4517p
L4 N3 N4 14.5699n
L5 N4 N5 68.6521n
L6 N5 N6 92.0413n
R1 2 N1 157.8926
R2 2 N2 25.8066
R3 2 N3 26.3545
R4 2 N4 26.6522
R5 2 N5 9.8403
R6 2 N6 8.5333
R7 2 N7 1.1054k
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760339A_3.9u 1 2
C1 1 N7 131.1918f
L1 1 N1 3.06u
L2 N1 N2 742.8370n
L3 N2 N3 819.2923p
L4 N3 N4 24.9908n
L5 N4 N5 84.3429n
L6 N5 N6 113.5388n
R1 2 N1 278.1925
R2 2 N2 26.9730
R3 2 N3 27.4690
R4 2 N4 27.9523
R5 2 N5 9.9662
R6 2 N6 8.6837
R7 2 N7 1.3709k
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760347A_4.7u 1 2
C1 1 N7 433.0876f
L1 1 N1 3.9977u
L2 N1 N2 734.0050n
L3 N2 N3 135.2855n
L4 N3 N4 72.2377n
L5 N4 N5 57.2282n
L6 N5 N6 287.7952n
R1 2 N1 198.1838
R2 2 N2 26.0714
R3 2 N3 26.9452
R4 2 N4 27.5069
R5 2 N5 9.8817
R6 2 N6 8.5409
R7 2 N7 784.6283
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760356A_5.6u 1 2
C1 1 N7 459.0344f
L1 1 N1 4.83u
L2 N1 N2 1.0405u
L3 N2 N3 816.1320p
L4 N3 N4 26.4147n
L5 N4 N5 13.1237n
L6 N5 N6 603.8984n
R1 2 N1 218.7445
R2 2 N2 25.3456
R3 2 N3 25.8975
R4 2 N4 26.2602
R5 2 N5 9.7824
R6 2 N6 8.5991
R7 2 N7 486.1824
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760382A_8.2u 1 2
C1 1 N7 291.6740f
L1 1 N1 7.3u
L2 N1 N2 1.2104u
L3 N2 N3 837.1269p
L4 N3 N4 91.4973n
L5 N4 N5 409.6341n
L6 N5 N6 1.3553u
R1 2 N1 272.5206
R2 2 N2 74.3932
R3 2 N3 54.3954
R4 2 N4 56.9118
R5 2 N5 16.4781
R6 2 N6 8.4993
R7 2 N7 851.0096
R8 2 1 10g
.ends 
*******
.subckt 0805A_744760410A_10u 1 2
C1 1 N7 204.4834f
L1 1 N1 8.9u
L2 N1 N2 1.7161u
L3 N2 N3 834.6607p
L4 N3 N4 77.5391n
L5 N4 N5 35.6154n
L6 N5 N6 9.7387u
R1 2 N1 481.9151
R2 2 N2 53.8234
R3 2 N3 53.8243
R4 2 N4 56.4302
R5 2 N5 10.9523
R6 2 N6 8.5315
R7 2 N7 1.1459k
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762312A_1.2u 1 2
C1 1 N7 158.7443f
L1 1 N1 1.15u
L2 N1 N2 25.7595n
L3 N2 N3 2.2471n
L4 N3 N4 35.0721n
L5 N4 N5 49.3056n
L6 N5 N6 26.2082n
R1 2 N1 37.0111
R2 2 N2 16.9448
R3 2 N3 20.1815
R4 2 N4 2.4163
R5 2 N5 9.4612
R6 2 N6 7.9902
R7 2 N7 171.5402
R8 2 1 10g
.ends 
******* 
.subckt 1008A_744762315A_1.5u 1 2
C1 1 N7 144.4482f
L1 1 N1 1.4750u
L2 N1 N2 43.4654n
L3 N2 N3 2.0276n
L4 N3 N4 43.3750n
L5 N4 N5 114.5311n
L6 N5 N6 51.8453n
R1 2 N1 39.7071
R2 2 N2 13.7898
R3 2 N3 18.0981
R4 2 N4 3.2315
R5 2 N5 9.4896
R6 2 N6 8.0124
R7 2 N7 138.0520
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762318A_1.8u 1 2
C1 1 N7 145.4549f
L1 1 N1 1.7850u
L2 N1 N2 57.9562n
L3 N2 N3 3.1587n
L4 N3 N4 9.8599n
L5 N4 N5 68.5705n
L6 N5 N6 27.6903n
R1 2 N1 34.3122
R2 2 N2 20.7754
R3 2 N3 23.0005
R4 2 N4 10.5653
R5 2 N5 9.5416
R6 2 N6 8.1049
R7 2 N7 109.6525
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762322A_2.2u 1 2
C1 1 N7 154.4785f
L1 1 N1 2.16u
L2 N1 N2 76.7015n
L3 N2 N3 4.5985n
L4 N3 N4 11.3131n
L5 N4 N5 72.6643n
L6 N5 N6 26.3276n
R1 2 N1 30.5560
R2 2 N2 21.9301
R3 2 N3 24.0282
R4 2 N4 15.3476
R5 2 N5 9.5424
R6 2 N6 8.1070
R7 2 N7 308.3232
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762327A_2.7u 1 2
C1 1 N7 377.6344f
L1 1 N1 2.65u
L2 N1 N2 120.7859n
L3 N2 N3 3.7238n
L4 N3 N4 7.2030n
L5 N4 N5 9.1192n
L6 N5 N6 4.6590n
R1 2 N1 24.5300
R2 2 N2 23.4744
R3 2 N3 29.1481
R4 2 N4 29.7704
R5 2 N5 20.5211
R6 2 N6 8.5261
R7 2 N7 172.7902
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762333A_3.3u 1 2
C1 1 N7 511.8368f
L1 1 N1 3.1u
L2 N1 N2 301.2330n
L3 N2 N3 744.1133p
L4 N3 N4 38.9127n
L5 N4 N5 47.9265n
L6 N5 N6 204.2512n
R1 2 N1 277.7959
R2 2 N2 26.2115
R3 2 N3 26.7451
R4 2 N4 27.1918
R5 2 N5 9.8920
R6 2 N6 8.5597
R7 2 N7 56.1459
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762339A_3.9u 1 2
C1 1 N7 713.2456f
L1 1 N1 3.6u
L2 N1 N2 182.3549n
L3 N2 N3 757.0463p
L4 N3 N4 139.0604n
L5 N4 N5 45.5489n
L6 N5 N6 2.0109u
R1 2 N1 142.0736
R2 2 N2 28.2253
R3 2 N3 28.6967
R4 2 N4 20.2129
R5 2 N5 9.9985
R6 2 N6 18.6399
R7 2 N7 135.2796
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762347A_4.7u 1 2
C1 1 N7 702.5978f
L1 1 N1 4.45u
L2 N1 N2 248.4266n
L3 N2 N3 757.2336p
L4 N3 N4 127.8327n
L5 N4 N5 51.0308n
L6 N5 N6 651.0043n
R1 2 N1 159.2400
R2 2 N2 28.7319
R3 2 N3 26.2849
R4 2 N4 25.4177
R5 2 N5 16.2226
R6 2 N6 19.2937
R7 2 N7 156.4933
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762356A_5.6u 1 2
C1 1 N7 323.8953f
L1 1 N1 5.1u
L2 N1 N2 605.4820n
L3 N2 N3 757.3560p
L4 N3 N4 327.1355n
L5 N4 N5 50.1316n
L6 N5 N6 588.7510n
R1 2 N1 185.5893
R2 2 N2 28.7002
R3 2 N3 26.2381
R4 2 N4 26.1783
R5 2 N5 18.6959
R6 2 N6 20.8881
R7 2 N7 268.1882
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762368A_6.8u 1 2
C1 1 N7 500.1575f
L1 1 N1 6.1u
L2 N1 N2 860.1723n
L3 N2 N3 761.1966p
L4 N3 N4 56.2783n
L5 N4 N5 59.2882n
L6 N5 N6 1.1711u
R1 2 N1 262.2656
R2 2 N2 30.7085
R3 2 N3 28.5802
R4 2 N4 28.9585
R5 2 N5 23.5813
R6 2 N6 21.3351
R7 2 N7 146.3916
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762382A_8.2u 1 2
C1 1 N7 730.0597f
L1 1 N1 7.25u
L2 N1 N2 962.4842n
L3 N2 N3 762.2250p
L4 N3 N4 60.3358n
L5 N4 N5 61.7402n
L6 N5 N6 2.2536u
R1 2 N1 265.8819
R2 2 N2 31.4736
R3 2 N3 29.4515
R4 2 N4 29.7693
R5 2 N5 24.4361
R6 2 N6 21.2667
R7 2 N7 127.7118
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762410A_10u 1 2
C1 1 N7 855.8897f
L1 1 N1 8.9u
L2 N1 N2 1.1434u
L3 N2 N3 762.6593p
L4 N3 N4 62.6732n
L5 N4 N5 63.2942n
L6 N5 N6 2.9201u
R1 2 N1 270.7618
R2 2 N2 32.1396
R3 2 N3 30.2058
R4 2 N4 30.4913
R5 2 N5 25.4603
R6 2 N6 21.1285
R7 2 N7 145.5541
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762415A_15u 1 2
C1 1 N7 365.0719f
L1 1 N1 14u
L2 N1 N2 2.6334u
L3 N2 N3 834.7144p
L4 N3 N4 77.5391n
L5 N4 N5 36.3963n
L6 N5 N6 9.8862u
R1 2 N1 558.8531
R2 2 N2 74.1014
R3 2 N3 64.1023
R4 2 N4 76.6831
R5 2 N5 21.3423
R6 2 N6 48.5308
R7 2 N7 109.0096
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762418A_18u 1 2
C1 1 N7 1.7966p
L1 1 N1 16.9u
L2 N1 N2 1.2439u
L3 N2 N3 836.0875p
L4 N3 N4 837.1967p
L5 N4 N5 269.6004n
L6 N5 N6 9.6504u
R1 2 N1 88.8571
R2 2 N2 55.2375
R3 2 N3 55.2405
R4 2 N4 25.7197
R5 2 N5 49.3684
R6 2 N6 18.5307
R7 2 N7 199.5243
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762422A_22u 1 2
C1 1 N7 564.1908f
L1 1 N1 20u
L2 N1 N2 2.2755u
L3 N2 N3 834.6409p
L4 N3 N4 834.7236p
L5 N4 N5 42.0581n
L6 N5 N6 1.2318u
R1 2 N1 339.4305
R2 2 N2 135.6962
R3 2 N3 133.7892
R4 2 N4 91.0732
R5 2 N5 36.1596
R6 2 N6 77.1113
R7 2 N7 264.3824
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762427A_27u 1 2
C1 1 N7 842.5091f
L1 1 N1 25u
L2 N1 N2 2.5507u
L3 N2 N3 835.3527p
L4 N3 N4 835.4006p
L5 N4 N5 42.3375n
L6 N5 N6 7.3808u
R1 2 N1 374.3260
R2 2 N2 259.8700
R3 2 N3 158.2613
R4 2 N4 130.9240
R5 2 N5 39.7641
R6 2 N6 126.2110
R7 2 N7 249.3839
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762433A_33u 1 2
C1 1 N7 887.1570f
L1 1 N1 30.3u
L2 N1 N2 3.1301u
L3 N2 N3 836.3149p
L4 N3 N4 836.3629p
L5 N4 N5 42.7424n
L6 N5 N6 7.6794u
R1 2 N1 371.5537
R2 2 N2 260.7929
R3 2 N3 160.6972
R4 2 N4 134.4474
R5 2 N5 40.1332
R6 2 N6 125.9908
R7 2 N7 228.6092
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762439A_39u 1 2
C1 1 N7 749.6654f
L1 1 N1 34.7u
L2 N1 N2 4.6998u
L3 N2 N3 835.9555p
L4 N3 N4 836.0075p
L5 N4 N5 43.6164n
L6 N5 N6 9.7186u
R1 2 N1 358.9162
R2 2 N2 267.3951
R3 2 N3 267.4135
R4 2 N4 177.2095
R5 2 N5 45.8166
R6 2 N6 127.5346
R7 2 N7 209.5201
R8 2 1 10g
.ends 
*******
.subckt 1008A_744762447A_47u 1 2
C1 1 N7 619.3667f
L1 1 N1 43.7u
L2 N1 N2 3.3960u
L3 N2 N3 836.2281p
L4 N3 N4 836.3151p
L5 N4 N5 46.4124n
L6 N5 N6 32.0350u
R1 2 N1 341.5274
R2 2 N2 294.2093
R3 2 N3 294.2254
R4 2 N4 235.2256
R5 2 N5 54.7054
R6 2 N6 129.2261
R7 2 N7 292.1897
R8 2 1 10g
.ends 
*******