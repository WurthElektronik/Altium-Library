**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  Toroidal PFC Chokes
* Matchcode:              WE-TORPFC
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Roberta    
* Date and Time:          2022-11-24
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com	
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt TOR37_760800401_118u 1 2
Rp 1 2 24.09k
Cp 1 2 4.21p
Rs 1 N3 14m
L1 N3 2 118u Rser = 0.00001
.ends TOR37_760800401_118u
*******
.subckt TOR37_760800403_355u 1 2
Rp 1 2 46.45k
Cp 1 2 7.71p
Rs 1 N3 27m
L1 N3 2 355u Rser = 0.00001
.ends TOR37_760800403_355u
*******
.subckt TOR37_760801401_118u 1 2
Rp 1 2 38.16k
Cp 1 2 3.81p
Rs 1 N3 14m
L1 N3 2 118u Rser = 0.00001
.ends TOR37_760801401_118u
*******
.subckt TOR37_760801403_355u 1 2
Rp 1 2 80.83k
Cp 1 2 6.82p
Rs 1 N3 27m
L1 N3 2 355u Rser = 0.00001
.ends TOR37_760801403_355u
*******
.subckt TOR50_760800201_194u 1 2
Rp 1 2 58.26k
Cp 1 2 4.98p
Rs 1 N3 27m
L1 N3 2 194u Rser = 0.00001
.ends TOR50_760800201_194u
*******
.subckt TOR50_760800202_389u 1 2
Rp 1 2 82.8k
Cp 1 2 7.38p
Rs 1 N3 37m
L1 N3 2 389u Rser = 0.00001
.ends TOR50_760800202_389u
*******
.subckt TOR50_760800203_584u 1 2
Rp 1 2 131.3k
Cp 1 2 12.07p
Rs 1 N3 53m
L1 N3 2 584u Rser = 0.00001
.ends TOR50_760800203_584u
*******
.subckt TOR50_760801201_194u 1 2
Rp 1 2 151.83k
Cp 1 2 3.46p
Rs 1 N3 27m
L1 N3 2 194u Rser = 0.00001
.ends TOR50_760801201_194u
*******
.subckt TOR50_760801202_389u 1 2
Rp 1 2 206.1k
Cp 1 2 6.81p
Rs 1 N3 37m
L1 N3 2 389u Rser = 0.00001
.ends TOR50_760801202_389u
*******
.subckt TOR50_760801203_584u 1 2
Rp 1 2 125k
Cp 1 2 11.1p
Rs 1 N3 53m
L1 N3 2 584u Rser = 0.00001
.ends TOR50_760801203_584u
*******
.subckt TOR43_760800101_255u 1 2
Rp 1 2 49.12k
Cp 1 2 4.69p
Rs 1 N3 28.8m
L1 N3 2 255u Rser = 0.00001
.ends TOR43_760800101_255u
*******
.subckt TOR43_760800102_510u 1 2
Rp 1 2 91.11k
Cp 1 2 5.15p
Rs 1 N3 44m
L1 N3 2 510u Rser = 0.00001
.ends TOR43_760800102_510u
*******
.subckt TOR43_760801101_255u 1 2
Rp 1 2 62.27k
Cp 1 2 2.57p
Rs 1 N3 29m
L1 N3 2 255u Rser = 0.00001
.ends TOR43_760801101_255u
*******
.subckt TOR43_760801102_510u 1 2
Rp 1 2 102.7k
Cp 1 2 4.04p
Rs 1 N3 44m
L1 N3 2 510u Rser = 0.00001
.ends TOR43_760801102_510u
*******
.subckt TOR75_760800301_180u 1 2
Rp 1 2 46.9k
Cp 1 2 11.58p
Rs 1 N3 18m
L1 N3 2 180u Rser = 0.00001
.ends TOR75_760800301_180u
*******
.subckt TOR75_760801301_180u 1 2
Rp 1 2 42.1k
Cp 1 2 11.84p
Rs 1 N3 18m
L1 N3 2 180u Rser = 0.00001
.ends TOR75_760801301_180u
*******
.subckt TOR75_760801321_720u 1 2
Rp 1 2 155k
Cp 1 2 6.27p
Rs 1 N3 34m
L1 N3 2 720u
.ends TOR75_760801321_720u
*******

