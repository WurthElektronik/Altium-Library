**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Resonant Converter
* Matchcode:              WE-LLCR
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Toby      
* Date and Time:          2022-05-17
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************

.subckt 760895751		12  10  15  14  1  5  3  7		
.param RxLkg=20624.15ohm					
.param Leakage=65uh					
Rlkg	12	12a	{RxLkg}		
L_Lkg	12	12a	{Leakage}	Rser=0.01mohm	
Lpri1	12a	10	335uH	Rser=64mohm	
Laux1	15	14	2.195uH	Rser=122mohm	
Lsec1	1	5	19.753uH	Rser=9.9mohm	
Lsec2	3	7	19.753uH	Rser=8.9mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=62.08pf					
.param Rdmp1=126917.83ohm					
Cpri1	12	10	{Cprm1}	Rser=10mohm	
Rdmp1	12	10	{Rdmp1}		
Rg3	12	0	20meg		
Rg5	15	0	20meg		
Rg7	10	0	20meg		
Rg9	14	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	5	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt 760895741		12  10  15  14  1  5  3  7		
.param RxLkg=23797.06ohm					
.param Leakage=65uh					
Rlkg	12	12a	{RxLkg}		
L_Lkg	12	12a	{Leakage}	Rser=0.01mohm	
Lpri1	12a	10	335uH	Rser=62.8mohm	
Laux1	15	14	2.195uH	Rser=124mohm	
Lsec1	1	5	4.938uH	Rser=3.6mohm	
Lsec2	3	7	4.938uH	Rser=4mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=46.63pf					
.param Rdmp1=146443.46ohm					
Cpri1	12	10	{Cprm1}	Rser=10mohm	
Rdmp1	12	10	{Rdmp1}		
Rg3	12	0	20meg		
Rg5	15	0	20meg		
Rg7	10	0	20meg		
Rg9	14	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	5	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt 760895731		12  10  15  14  1  5  3  7		
.param RxLkg=30336.48ohm					
.param Leakage=100uh					
Rlkg	12	12a	{RxLkg}		
L_Lkg	12	12a	{Leakage}	Rser=0.01mohm	
Lpri1	12a	10	375uH	Rser=106mohm	
Laux1	15	14	3.49uH	Rser=150mohm	
Lsec1	1	5	1.551uH	Rser=2.7mohm	
Lsec2	3	7	1.551uH	Rser=2.9mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=57.19pf					
.param Rdmp1=144098.26ohm					
Cpri1	12	10	{Cprm1}	Rser=10mohm	
Rdmp1	12	10	{Rdmp1}		
Rg3	12	0	20meg		
Rg5	15	0	20meg		
Rg7	10	0	20meg		
Rg9	14	0	20meg		
Rg11	1	0	20meg		
Rg12	3	0	20meg		
Rg19	5	0	20meg		
Rg20	7	0	20meg		
.ends					

.subckt 760895651		4  2  5  6  8  12  10  14		
.param RxLkg=29204.06ohm					
.param Leakage=95uh					
Rlkg	4	4a	{RxLkg}		
L_Lkg	4	4a	{Leakage}	Rser=0.01mohm	
Lpri1	4a	2	405uH	Rser=121mohm	
Laux1	5	6	3.673uH	Rser=139mohm	
Lsec1	8	12	26.122uH	Rser=17.9mohm	
Lsec2	10	14	26.122uH	Rser=17.9mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=52.91pf					
.param Rdmp1=153705.56ohm					
Cpri1	4	2	{Cprm1}	Rser=10mohm	
Rdmp1	4	2	{Rdmp1}		
Rg3	4	0	20meg		
Rg5	5	0	20meg		
Rg7	2	0	20meg		
Rg9	6	0	20meg		
Rg11	8	0	20meg		
Rg12	10	0	20meg		
Rg19	12	0	20meg		
Rg20	14	0	20meg		
.ends					

.subckt 760895641		4  2  5  6  8  12  10  14		
.param RxLkg=26605.14ohm					
.param Leakage=95uh					
Rlkg	4	4a	{RxLkg}		
L_Lkg	4	4a	{Leakage}	Rser=0.01mohm	
Lpri1	4a	2	405uH	Rser=120mohm	
Laux1	5	6	3.673uH	Rser=137mohm	
Lsec1	8	12	6.531uH	Rser=6.4mohm	
Lsec2	10	14	6.531uH	Rser=6.3mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=63.75pf					
.param Rdmp1=140027.07ohm					
Cpri1	4	2	{Cprm1}	Rser=10mohm	
Rdmp1	4	2	{Rdmp1}		
Rg3	4	0	20meg		
Rg5	5	0	20meg		
Rg7	2	0	20meg		
Rg9	6	0	20meg		
Rg11	8	0	20meg		
Rg12	10	0	20meg		
Rg19	12	0	20meg		
Rg20	14	0	20meg		
.ends					

.subckt 760895631		4  2  5  6  8  11  10  13		
.param RxLkg=30080.91ohm					
.param Leakage=95uh					
Rlkg	4	4a	{RxLkg}		
L_Lkg	4	4a	{Leakage}	Rser=0.01mohm	
Lpri1	4a	2	405uH	Rser=123mohm	
Laux1	5	6	3.673uH	Rser=128mohm	
Lsec1	8	11	1.633uH	Rser=2.2mohm	
Lsec2	10	13	1.633uH	Rser=2mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=49.87pf					
.param Rdmp1=158320.56ohm					
Cpri1	4	2	{Cprm1}	Rser=10mohm	
Rdmp1	4	2	{Rdmp1}		
Rg3	4	0	20meg		
Rg5	5	0	20meg		
Rg7	2	0	20meg		
Rg9	6	0	20meg		
Rg11	8	0	20meg		
Rg12	10	0	20meg		
Rg19	11	0	20meg		
Rg20	13	0	20meg		
.ends					

.subckt 760895451		4  2  5  6  8  10  9  11		
.param RxLkg=29850.79ohm					
.param Leakage=100uh					
Rlkg	4	4a	{RxLkg}		
L_Lkg	4	4a	{Leakage}	Rser=0.01mohm	
Lpri1	4a	2	500uH	Rser=228.5mohm	
Laux1	5	6	4.408uH	Rser=128mohm	
Lsec1	8	10	31.347uH	Rser=22.8mohm	
Lsec2	9	11	31.347uH	Rser=22.9mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=46.76pf					
.param Rdmp1=179104.71ohm					
Cpri1	4	2	{Cprm1}	Rser=10mohm	
Rdmp1	4	2	{Rdmp1}		
Rg3	4	0	20meg		
Rg5	5	0	20meg		
Rg7	2	0	20meg		
Rg9	6	0	20meg		
Rg11	8	0	20meg		
Rg12	9	0	20meg		
Rg19	10	0	20meg		
Rg20	11	0	20meg		
.ends					

.subckt 760895441		4  2  5  6  8  10  9  11		
.param RxLkg=32592.14ohm					
.param Leakage=100uh					
Rlkg	4	4a	{RxLkg}		
L_Lkg	4	4a	{Leakage}	Rser=0.01mohm	
Lpri1	4a	2	500uH	Rser=237mohm	
Laux1	5	6	4.408uH	Rser=121.7mohm	
Lsec1	8	10	7.837uH	Rser=7.4mohm	
Lsec2	9	11	7.837uH	Rser=7.4mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=39.225pf					
.param Rdmp1=195552.83ohm					
Cpri1	4	2	{Cprm1}	Rser=10mohm	
Rdmp1	4	2	{Rdmp1}		
Rg3	4	0	20meg		
Rg5	5	0	20meg		
Rg7	2	0	20meg		
Rg9	6	0	20meg		
Rg11	8	0	20meg		
Rg12	9	0	20meg		
Rg19	10	0	20meg		
Rg20	11	0	20meg		
.ends					

.subckt 760895431		4  2  5  6  8  10  9  11		
.param RxLkg=31739.51ohm					
.param Leakage=100uh					
Rlkg	4	4a	{RxLkg}		
L_Lkg	4	4a	{Leakage}	Rser=0.01mohm	
Lpri1	4a	2	500uH	Rser=229mohm	
Laux1	5	6	4.408uH	Rser=121.7mohm	
Lsec1	8	10	1.959uH	Rser=2.88mohm	
Lsec2	9	11	1.959uH	Rser=2.3mohm	
K Lpri1  Laux1  Lsec1 Lsec2       1					
.param Cprm1=41.36pf					
.param Rdmp1=190437.06ohm					
Cpri1	4	2	{Cprm1}	Rser=10mohm	
Rdmp1	4	2	{Rdmp1}		
Rg3	4	0	20meg		
Rg5	5	0	20meg		
Rg7	2	0	20meg		
Rg9	6	0	20meg		
Rg11	8	0	20meg		
Rg12	9	0	20meg		
Rg19	10	0	20meg		
Rg20	11	0	20meg		
.ends					
