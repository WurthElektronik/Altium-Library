**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  MLCCs - Multilayer Ceramic Chip Capacitors
* Matchcode:              WCAP-CSMH
* Library Type:           spice
* Version:                rev
* Created/modified by:    Ella
* Date and Time:          5/20/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0603_885342006001_10pF 1 2
Rser 1 3 0.526591507248
Lser 2 4 6.5841246E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885342006001_10pF
*******
.subckt 0603_885342006002_33pF 1 2
Rser 1 3 0.255116824504
Lser 2 4 5.30449805E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885342006002_33pF
*******
.subckt 0603_885342006003_100pF 1 2
Rser 1 3 0.146495221684
Lser 2 4 4.78406333E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885342006003_100pF
*******
.subckt 0603_885342206001_100pF 1 2
Rser 1 3 0.897508199816
Lser 2 4 3.40719264E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885342206001_100pF
*******
.subckt 0603_885342006004_220pF 1 2
Rser 1 3 0.0871099668085
Lser 2 4 4.10447243E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885342006004_220pF
*******
.subckt 0603_885342206002_330pF 1 2
Rser 1 3 0.459205969757
Lser 2 4 3.62972471E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885342206002_330pF
*******
.subckt 0603_885342006005_470pF 1 2
Rser 1 3 0.0832834441759
Lser 2 4 4.18832836E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885342006005_470pF
*******
.subckt 0603_885342206003_1nF 1 2
Rser 1 3 0.229494082774
Lser 2 4 4.2835564E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885342206003_1nF
*******
.subckt 0603_885342206004_1.5nF 1 2
Rser 1 3 0.178697894647
Lser 2 4 3.79706604E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885342206004_1.5nF
*******
.subckt 0603_885342206005_3.3nF 1 2
Rser 1 3 0.147147912937
Lser 2 4 3.75939961E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885342206005_3.3nF
*******
.subckt 0603_885342206006_10nF 1 2
Rser 1 3 0.056712206124
Lser 2 4 4.04185706E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885342206006_10nF
*******
.subckt 0805_885342007004_15pF 1 2
Rser 1 3 0.213471971511
Lser 2 4 4.77553318E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885342007004_15pF
*******
.subckt 0805_885342007006_47pF 1 2
Rser 1 3 0.146554502609
Lser 2 4 4.81671007E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885342007006_47pF
*******
.subckt 0805_885342207001_100pF 1 2
Rser 1 3 0.132042743101
Lser 2 4 3.82973241E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885342207001_100pF
*******
.subckt 0805_885342207015_100pF 1 2
Rser 1 3 1.46345969291
Lser 2 4 4.01548958E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885342207015_100pF
*******
.subckt 0805_885342007001_220pF 1 2
Rser 1 3 0.0850728682842
Lser 2 4 3.94126801E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885342007001_220pF
*******
.subckt 0805_885342007002_330pF 1 2
Rser 1 3 0.062685416378
Lser 2 4 4.11124644E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885342007002_330pF
*******
.subckt 0805_885342207002_470pF 1 2
Rser 1 3 0.189434542942
Lser 2 4 3.77514445E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885342207002_470pF
*******
.subckt 0805_885342207007_470pF 1 2
Rser 1 3 0.963404301108
Lser 2 4 4.41658976E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885342207007_470pF
*******
.subckt 0805_885342207012_470pF 1 2
Rser 1 3 0.0118150527569
Lser 2 4 4.45623546E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885342207012_470pF
*******
.subckt 0805_885342007003_1nF 1 2
Rser 1 3 0.0804888218968
Lser 2 4 4.05575252E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885342007003_1nF
*******
.subckt 0805_885342207003_1nF 1 2
Rser 1 3 0.217753942776
Lser 2 4 4.3508637E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885342207003_1nF
*******
.subckt 0805_885342207008_1nF 1 2
Rser 1 3 0.258021361158
Lser 2 4 4.18753287E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885342207008_1nF
*******
.subckt 0805_885342207013_1nF 1 2
Rser 1 3 0.275047233421
Lser 2 4 4.12151413E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885342207013_1nF
*******
.subckt 0805_885342007005_2.2nF 1 2
Rser 1 3 0.0664836922917
Lser 2 4 2.47874891E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885342007005_2.2nF
*******
.subckt 0805_885342207016_2.2nF 1 2
Rser 1 3 0.0818041012502
Lser 2 4 3.76209238E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885342207016_2.2nF
*******
.subckt 0805_885342207004_4.7nF 1 2
Rser 1 3 0.107
Lser 2 4 0.0000000009
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885342207004_4.7nF
*******
.subckt 0805_885342207009_4.7nF 1 2
Rser 1 3 0.394840579191
Lser 2 4 4.45623453E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885342207009_4.7nF
*******
.subckt 0805_885342207005_10nF 1 2
Rser 1 3 0.07
Lser 2 4 0.0000000011
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885342207005_10nF
*******
.subckt 0805_885342207010_10nF 1 2
Rser 1 3 0.0485521865845
Lser 2 4 4.34329744E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885342207010_10nF
*******
.subckt 0805_885342207014_10nF 1 2
Rser 1 3 0.0478133926287
Lser 2 4 3.58284831E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885342207014_10nF
*******
.subckt 0805_885342207006_22nF 1 2
Rser 1 3 0.0324448031493
Lser 2 4 3.75007753E-10
C1 3 4 0.000000022
Rpar 3 4 4540000000
.ends 0805_885342207006_22nF
*******
.subckt 0805_885342207011_22nF 1 2
Rser 1 3 0.0345951343679
Lser 2 4 3.77731639E-10
C1 3 4 0.000000022
Rpar 3 4 4540000000
.ends 0805_885342207011_22nF
*******
.subckt 1206_885342008008_22pF 1 2
Rser 1 3 0.209638135659
Lser 2 4 5.17238769E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1206_885342008008_22pF
*******
.subckt 1206_885342008001_47pF 1 2
Rser 1 3 0.197952268363
Lser 2 4 5.47249965E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885342008001_47pF
*******
.subckt 1206_885342008010_68pF 1 2
Rser 1 3 0.118896244952
Lser 2 4 5.50065477E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 1206_885342008010_68pF
*******
.subckt 1206_885342008004_100pF 1 2
Rser 1 3 0.135674317711
Lser 2 4 4.77445122E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885342008004_100pF
*******
.subckt 1206_885342008009_100pF 1 2
Rser 1 3 0.103584713826
Lser 2 4 5.23151691E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885342008009_100pF
*******
.subckt 1206_885342008011_100pF 1 2
Rser 1 3 0.0971330396442
Lser 2 4 4.9235317E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885342008011_100pF
*******
.subckt 1206_885342208022_100pF 1 2
Rser 1 3 0.753874561624
Lser 2 4 1.96091472E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885342208022_100pF
*******
.subckt 1206_885342208016_150pF 1 2
Rser 1 3 0.685541200809
Lser 2 4 4.45467633E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885342208016_150pF
*******
.subckt 1206_885342008002_220pF 1 2
Rser 1 3 0.0989171163333
Lser 2 4 4.16981088E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885342008002_220pF
*******
.subckt 1206_885342208005_470pF 1 2
Rser 1 3 0.385869412824
Lser 2 4 5.28105714E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885342208005_470pF
*******
.subckt 1206_885342208017_470pF 1 2
Rser 1 3 0.436768993856
Lser 2 4 6.28786815E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885342208017_470pF
*******
.subckt 1206_885342208023_470pF 1 2
Rser 1 3 0.39020934864
Lser 2 4 5.13086603E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885342208023_470pF
*******
.subckt 1206_885342008003_1nF 1 2
Rser 1 3 0.0609307626631
Lser 2 4 4.05708124E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885342008003_1nF
*******
.subckt 1206_885342008005_1nF 1 2
Rser 1 3 0.0380244845246
Lser 2 4 2.9643754E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885342008005_1nF
*******
.subckt 1206_885342208006_1nF 1 2
Rser 1 3 0.177597971676
Lser 2 4 4.56580055E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885342208006_1nF
*******
.subckt 1206_885342208011_1nF 1 2
Rser 1 3 0.192424270317
Lser 2 4 4.48778059E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885342208011_1nF
*******
.subckt 1206_885342208018_1nF 1 2
Rser 1 3 0.22866226126
Lser 2 4 4.63515197E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885342208018_1nF
*******
.subckt 1206_885342208024_1nF 1 2
Rser 1 3 0.147813230311
Lser 2 4 1.64762577E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885342208024_1nF
*******
.subckt 1206_885342008006_1.5nF 1 2
Rser 1 3 0.0298853431351
Lser 2 4 3.033024E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885342008006_1.5nF
*******
.subckt 1206_885342008007_2.2nF 1 2
Rser 1 3 0.0317456317923
Lser 2 4 6.20552358E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885342008007_2.2nF
*******
.subckt 1206_885342208007_2.2nF 1 2
Rser 1 3 0.144882392111
Lser 2 4 4.63500612E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885342208007_2.2nF
*******
.subckt 1206_885342208019_2.2nF 1 2
Rser 1 3 0.15123586699
Lser 2 4 4.79802798E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885342208019_2.2nF
*******
.subckt 1206_885342208008_4.7nF 1 2
Rser 1 3 0.0789077852137
Lser 2 4 4.84745669E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885342208008_4.7nF
*******
.subckt 1206_885342208020_4.7nF 1 2
Rser 1 3 0.0932877077493
Lser 2 4 4.87623506E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885342208020_4.7nF
*******
.subckt 1206_885342208003_10nF 1 2
Rser 1 3 0.098296958648
Lser 2 4 4.63188389E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885342208003_10nF
*******
.subckt 1206_885342208009_10nF 1 2
Rser 1 3 0.0970703444071
Lser 2 4 4.20580769E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885342208009_10nF
*******
.subckt 1206_885342208012_10nF 1 2
Rser 1 3 0.0892072672408
Lser 2 4 4.20340712E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885342208012_10nF
*******
.subckt 1206_885342208021_10nF 1 2
Rser 1 3 0.0745593249743
Lser 2 4 1.289927921E-09
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885342208021_10nF
*******
.subckt 1206_885342208013_15nF 1 2
Rser 1 3 0.0419773550564
Lser 2 4 5.14619153E-10
C1 3 4 0.000000015
Rpar 3 4 6660000000
.ends 1206_885342208013_15nF
*******
.subckt 1206_885342208001_22nF 1 2
Rser 1 3 0.106950110433
Lser 2 4 7.34881047E-10
C1 3 4 0.000000022
Rpar 3 4 4540000000
.ends 1206_885342208001_22nF
*******
.subckt 1206_885342208010_22nF 1 2
Rser 1 3 0.0723894054808
Lser 2 4 5.26703102E-10
C1 3 4 0.000000022
Rpar 3 4 4540000000
.ends 1206_885342208010_22nF
*******
.subckt 1206_885342208014_22nF 1 2
Rser 1 3 0.0616439765027
Lser 2 4 4.76808143E-10
C1 3 4 0.000000022
Rpar 3 4 4540000000
.ends 1206_885342208014_22nF
*******
.subckt 1206_885342208015_33nF 1 2
Rser 1 3 0.0550803748741
Lser 2 4 5.09753727E-10
C1 3 4 0.000000033
Rpar 3 4 3030000000
.ends 1206_885342208015_33nF
*******
.subckt 1206_885342208026_47nF 1 2
Rser 1 3 0.025
Lser 2 4 0.00000000093
C1 3 4 0.000000047
Rpar 3 4 2127000000
.ends 1206_885342208026_47nF
*******
.subckt 1206_885342208002_100nF 1 2
Rser 1 3 0.0312255702324
Lser 2 4 4.59358937E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1206_885342208002_100nF
*******
.subckt 1206_885342208004_100nF 1 2
Rser 1 3 0.023410869744
Lser 2 4 6.25812228E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1206_885342208004_100nF
*******
.subckt 1210_885342009004_10pF 1 2
Rser 1 3 0.259686916806
Lser 2 4 3.16360399E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1210_885342009004_10pF
*******
.subckt 1210_885342009002_22pF 1 2
Rser 1 3 0.229015378654
Lser 2 4 2.60728331E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1210_885342009002_22pF
*******
.subckt 1210_885342009005_220pF 1 2
Rser 1 3 0.110218233392
Lser 2 4 3.96893935E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1210_885342009005_220pF
*******
.subckt 1210_885342209008_220pF 1 2
Rser 1 3 0.480745779266
Lser 2 4 3.58505408E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1210_885342209008_220pF
*******
.subckt 1210_885342009003_1nF 1 2
Rser 1 3 0.0569267068127
Lser 2 4 3.92362421E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885342009003_1nF
*******
.subckt 1210_885342209006_1nF 1 2
Rser 1 3 0.194650555528
Lser 2 4 3.7524441E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885342209006_1nF
*******
.subckt 1210_885342209009_1nF 1 2
Rser 1 3 0.343504568556
Lser 2 4 3.91503622E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885342209009_1nF
*******
.subckt 1210_885342009001_4.7nF 1 2
Rser 1 3 0.0281181269798
Lser 2 4 3.85364184E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1210_885342009001_4.7nF
*******
.subckt 1210_885342009007_5.6nF 1 2
Rser 1 3 0.0198
Lser 2 4 0.00000000065
C1 3 4 0.0000000056
Rpar 3 4 10000000000
.ends 1210_885342009007_5.6nF
*******
.subckt 1210_885342209001_15nF 1 2
Rser 1 3 0.0483587105706
Lser 2 4 2.82691432E-10
C1 3 4 0.000000015
Rpar 3 4 6660000000
.ends 1210_885342209001_15nF
*******
.subckt 1210_885342209007_22nF 1 2
Rser 1 3 0.0235915106864
Lser 2 4 3.40725306E-10
C1 3 4 0.000000022
Rpar 3 4 4550000000
.ends 1210_885342209007_22nF
*******
.subckt 1210_885342209004_33nF 1 2
Rser 1 3 0.0267458879248
Lser 2 4 3.56097176E-10
C1 3 4 0.000000033
Rpar 3 4 3030000000
.ends 1210_885342209004_33nF
*******
.subckt 1210_885342209005_68nF 1 2
Rser 1 3 0.0142659341117
Lser 2 4 4.38758468E-10
C1 3 4 0.000000068
Rpar 3 4 1470000000
.ends 1210_885342209005_68nF
*******
.subckt 1210_885342209002_100nF 1 2
Rser 1 3 0.0176148022492
Lser 2 4 6.26675864E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1210_885342209002_100nF
*******
.subckt 1210_885342209003_220nF 1 2
Rser 1 3 0.0155
Lser 2 4 0.00000000109
C1 3 4 0.00000022
Rpar 3 4 450000000
.ends 1210_885342209003_220nF
*******
.subckt 1808_885342010001_10pF 1 2
Rser 1 3 0.383139788341
Lser 2 4 6.2563052E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1808_885342010001_10pF
*******
.subckt 1808_885342010002_68pF 1 2
Rser 1 3 0.199225923302
Lser 2 4 6.41922587E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 1808_885342010002_68pF
*******
.subckt 1808_885342010003_100pF 1 2
Rser 1 3 0.187678931908
Lser 2 4 3.95010123E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1808_885342010003_100pF
*******
.subckt 1808_885342210003_470pF 1 2
Rser 1 3 0.249636437656
Lser 2 4 6.86223834E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1808_885342210003_470pF
*******
.subckt 1808_885342210001_1nF 1 2
Rser 1 3 0.251539206056
Lser 2 4 0.000000000675676
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1808_885342210001_1nF
*******
.subckt 1808_885342210004_1nF 1 2
Rser 1 3 0.266638508594
Lser 2 4 5.71850465E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1808_885342210004_1nF
*******
.subckt 1808_885342210002_2.2nF 1 2
Rser 1 3 0.155849577263
Lser 2 4 1.020120375E-09
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1808_885342210002_2.2nF
*******
.subckt 1812_885342011002_100pF 1 2
Rser 1 3 0.189291210432
Lser 2 4 5.09926281E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1812_885342011002_100pF
*******
.subckt 1812_885342011001_1nF 1 2
Rser 1 3 0.0857100266727
Lser 2 4 5.61273281E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_885342011001_1nF
*******
.subckt 1812_885342211009_1nF 1 2
Rser 1 3 0.24385903253
Lser 2 4 5.78618732E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_885342211009_1nF
*******
.subckt 1812_885342011003_1.5nF 1 2
Rser 1 3 0.0341746658869
Lser 2 4 7.61664077E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1812_885342011003_1.5nF
*******
.subckt 1812_885342211007_2.2nF 1 2
Rser 1 3 0.0585952173592
Lser 2 4 3.85402312E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1812_885342211007_2.2nF
*******
.subckt 1812_885342211010_2.2nF 1 2
Rser 1 3 0.133897819821
Lser 2 4 5.96006665E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1812_885342211010_2.2nF
*******
.subckt 1812_885342211001_4.7nF 1 2
Rser 1 3 0.0023387168803
Lser 2 4 1.249851605E-09
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1812_885342211001_4.7nF
*******
.subckt 1812_885342211008_4.7nF 1 2
Rser 1 3 0.157731534341
Lser 2 4 5.5102414E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1812_885342211008_4.7nF
*******
.subckt 1812_885342211004_10nF 1 2
Rser 1 3 0.0909203279595
Lser 2 4 3.1100596E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885342211004_10nF
*******
.subckt 1812_885342211002_100nF 1 2
Rser 1 3 0.0217199364802
Lser 2 4 6.76406598E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1812_885342211002_100nF
*******
.subckt 1812_885342211005_100nF 1 2
Rser 1 3 0.0140466361405
Lser 2 4 8.57894111E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1812_885342211005_100nF
*******
.subckt 1812_885342211006_100nF 1 2
Rser 1 3 0.0138355219015
Lser 2 4 8.12989182E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1812_885342211006_100nF
*******
.subckt 1812_885342211003_470nF 1 2
Rser 1 3 0.00691642348128
Lser 2 4 8.54557411E-10
C1 3 4 0.00000047
Rpar 3 4 210000000
.ends 1812_885342211003_470nF
*******
.subckt 2220_885342014230_100pF 1 2
Rser 1 3 0.14
Lser 2 4 0.0000000011
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 2220_885342014230_100pF
*******
.subckt 2220_885342214216_22nF 1 2
Rser 1 3 0.0350214797086
Lser 2 4 1.242206564E-09
C1 3 4 0.000000022
Rpar 3 4 5000000000
.ends 2220_885342214216_22nF
*******
.subckt 2220_885342214173_100nF 1 2
Rser 1 3 0.0165
Lser 2 4 0.000000001
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 2220_885342214173_100nF
*******
.subckt 2220_885342214142_220nF 1 2
Rser 1 3 0.0165
Lser 2 4 0.000000001
C1 3 4 0.00000022
Rpar 3 4 500000000
.ends 2220_885342214142_220nF
*******
.subckt 2220_885342214001_1uF 1 2
Rser 1 3 0.0064
Lser 2 4 0.0000000013
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 2220_885342214001_1uF
*******
.subckt 2220_885342214002_1uF 1 2
Rser 1 3 0.0084
Lser 2 4 0.0000000011
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 2220_885342214002_1uF
*******
.subckt 2220_885342214003_2.2uF 1 2
Rser 1 3 0.0053
Lser 2 4 0.000000001
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 2220_885342214003_2.2uF
*******
