**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Full-color Chip LED Diffused
* Matchcode:              WL-SFCD
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-16
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0606_150066M153000 1 2 3 4
D1 4 1 Red
.MODEL Red D
+ IS=10.000E-21
+ N=1.7618
+ RS=1.0000E-6
+ IKF=2.0622E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D2 4 2 Green
.MODEL Green D
+ IS=9.0185E-15
+ N=4.0502
+ RS=.65833
+ IKF=796.05E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D3 4 3 Blue
.MODEL Blue D
+ IS=13.286E-15
+ N=4.2265
+ RS=.69984
+ IKF=801.48E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
****************************
.subckt 0805_150080M153000 1 2 3 4
D1 4 1 Red
.MODEL Red D
+ IS=10.000E-21
+ N=1.7618
+ RS=1.0000E-6
+ IKF=2.0622E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D2 4 2 Green
.MODEL Green D
+ IS=24.280E-12
+ N=3.8516
+ RS=1.1745
+ IKF=792.64E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D3 4 3 Blue
.MODEL Blue D
+ IS=847.93E-18
+ N=3.4400
+ RS=.51865
+ IKF=753.31E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
****************************
.subckt 1210_150121M153000 1 2 3 4
D1 4 1 Red
.MODEL Red D
+ IS=10.000E-21
+ N=1.7618
+ RS=1.0000E-6
+ IKF=2.0622E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D2 4 2 Green
.MODEL Green D
+ IS=847.93E-18
+ N=3.4400
+ RS=.51865
+ IKF=753.31E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
D3 4 3 Blue
.MODEL Blue D
+ IS=24.280E-12
+ N=3.8516
+ RS=1.1745
+ IKF=792.64E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
************************