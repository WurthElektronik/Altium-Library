**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  EMI Multilayer Power Suppression Bead
* Matchcode:              WE-MPSA 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-30
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0805_78279220321_320Ohm 1 2
Rp 1 2 346.395
Cp 1 2 .917706p
L1 N3 2 .977736u
Rs 1 N3 .05
.ends 0805_78279220321_320Ohm
*******
.subckt 0805_78279220601_600Ohm 1 2
Rp 1 2 551.262
Cp 1 2 1.201p
L1 N3 2 1.803u
Rs 1 N3 .08
.ends 0805_78279220601_600Ohm
*******
.subckt 0805_78279220800_80Ohm 1 2
Rp 1 2 118.851
Cp 1 2 .250382p
L1 N3 2 .23556u
Rs 1 N3 .018
.ends 0805_78279220800_80Ohm
*******
.subckt 1206_78279221281_280Ohm 1 2
Rp 1 2 286.254
Cp 1 2 2.056p
L1 N3 2 .82817u
Rs 1 N3 .035
.ends 1206_78279221281_280Ohm
*******
.subckt 1206_78279221601_600Ohm 1 2
Rp 1 2 606.641
Cp 1 2 2.114p
L1 N3 2 1.793u
Rs 1 N3 .05
.ends 1206_78279221601_600Ohm
*******
.subckt 1612_78279223560_56Ohm 1 2
Rp 1 2 88.557
Cp 1 2 .175113p
L1 N3 2 .139605u
Rs 1 N3 .004
.ends 1612_78279223560_56Ohm
*******
.subckt 2220_78279224101_100Ohm 1 2
Rp 1 2 158.28
Cp 1 2 .099884p
L1 N3 2 .244751u
Rs 1 N3 .005
.ends 2220_78279224101_100Ohm
*******
.subckt 2220_78279224151_150Ohm 1 2
Rp 1 2 229.326
Cp 1 2 .135469p
L1 N3 2 .401877u
Rs 1 N3 .01
.ends 2220_78279224151_150Ohm
*******
.subckt 2220_78279224171_170Ohm 1 2
Rp 1 2 282.509
Cp 1 2 .106992p
L1 N3 2 .433549u
Rs 1 N3 .015
.ends 2220_78279224171_170Ohm
*******
.subckt 2220_78279224181_180Ohm 1 2
Rp 1 2 239.53
Cp 1 2 .140769p
L1 N3 2 .491744u
Rs 1 N3 .01
.ends 2220_78279224181_180Ohm
*******
.subckt 2220_78279224251_250Ohm 1 2
Rp 1 2 302.04
Cp 1 2 1.257p
L1 N3 2 .837627u
Rs 1 N3 .012
.ends 2220_78279224251_250Ohm
*******
.subckt 2220_78279224271_270Ohm 1 2
Rp 1 2 353.295
Cp 1 2 .339305p
L1 N3 2 .933918u
Rs 1 N3 .02
.ends 2220_78279224271_270Ohm
*******
.subckt 2220_78279224401_400Ohm 1 2
Rp 1 2 463.919
Cp 1 2 1.486p
L1 N3 2 1.578u
Rs 1 N3 .02
.ends 2220_78279224401_400Ohm
*******
.subckt 2220_78279224551_550Ohm 1 2
Rp 1 2 665.899
Cp 1 2 .231507p
L1 N3 2 1.369u
Rs 1 N3 .035
.ends 2220_78279224551_550Ohm
*******
.subckt 3312_78279225101_100Ohm 1 2
Rp 1 2 160.523
Cp 1 2 .059432p
L1 N3 2 .275642u
Rs 1 N3 .004
.ends 3312_78279225101_100Ohm
*******
.subckt 1812_78279226101_100Ohm 1 2
Rp 1 2 157.085
Cp 1 2 .087376p
L1 N3 2 .238388u
Rs 1 N3 .006
.ends 1812_78279226101_100Ohm
*******
