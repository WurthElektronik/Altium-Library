**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Multilayer Ceramic SMT Inductor 
* Matchcode:              WE-MK 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-24
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0201_7447820010_1n 1 2
C1 1 N7 252.6464f
L1 1 N1 0.95n
L2 N1 N2 219.3834p
L3 N2 N3 343.0117p
L4 N3 N4 459.3208p
L5 N4 N5 77.2700p
L6 N5 N6 54.4817p
R1 2 N1 453.2257m
R2 2 N2 197.3924m
R3 2 N3 434.9411m
R4 2 N4 392.5233m
R5 2 N5 348.7678m
R6 2 N6 96.5857m
R7 2 N7 1.9655
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820012_1.2n 1 2
C1 1 N7 0.2p
L1 1 N1 1.15n
L2 N1 N2 247.8759p
L3 N2 N3 343.7710p
L4 N3 N4 460.0589p
L5 N4 N5 77.2770p
L6 N5 N6 54.4873p
R1 2 N1 530.8745m
R2 2 N2 199.8839m
R3 2 N3 435.5468m
R4 2 N4 393.2090m
R5 2 N5 349.5902m
R6 2 N6 96.6861m
R7 2 N7 1.9668
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820015_1.5n 1 2
C1 1 N7 0.15p
L1 1 N1 1.3n
L2 N1 N2 200.4664p
L3 N2 N3 399.6617p
L4 N3 N4 495.4626p
L5 N4 N5 77.5313p
L6 N5 N6 54.6490p
R1 2 N1 719.2764m
R2 2 N2 344.4866m
R3 2 N3 456.1688m
R4 2 N4 402.5555m
R5 2 N5 359.0284m
R6 2 N6 97.7494m
R7 2 N7 1.9706
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820018_1.8n 1 2
C1 1 N7 0.14p
L1 1 N1 1.7n
L2 N1 N2 335.7177p
L3 N2 N3 596.4608p
L4 N3 N4 706.6429p
L5 N4 N5 79.1069p
L6 N5 N6 55.6649p
R1 2 N1 825.9598m
R2 2 N2 317.3420m
R3 2 N3 532.8549m
R4 2 N4 460.9317m
R5 2 N5 418.9950m
R6 2 N6 105.2425m
R7 2 N7 1.9764
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820020_2n 1 2
C1 1 N7 0.16p
L1 1 N1 1.8n
L2 N1 N2 201.6446p
L3 N2 N3 623.6153p
L4 N3 N4 747.7181p
L5 N4 N5 79.4118p
L6 N5 N6 55.8564p
R1 2 N1 593.6751m
R2 2 N2 205.9029m
R3 2 N3 540.5001m
R4 2 N4 473.3010m
R5 2 N5 431.9246m
R6 2 N6 107.1230m
R7 2 N7 1.9727
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820022_2.2n 1 2
C1 1 N7 0.14p
L1 1 N1 2n
L2 N1 N2 364.2086p
L3 N2 N3 637.5231p
L4 N3 N4 755.6190p
L5 N4 N5 79.4712p
L6 N5 N6 55.8973p
R1 2 N1 742.9116m
R2 2 N2 300.6071m
R3 2 N3 545.9497m
R4 2 N4 474.8793m
R5 2 N5 433.3975m
R6 2 N6 107.3178m
R7 2 N7 1.9758
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820024_2.4n 1 2
C1 1 N7 0.15p
L1 1 N1 2.2n
L2 N1 N2 379.9885p
L3 N2 N3 637.0462p
L4 N3 N4 755.3142p
L5 N4 N5 79.4707p
L6 N5 N6 55.8982p
R1 2 N1 787.4117m
R2 2 N2 299.8665m
R3 2 N3 545.7213m
R4 2 N4 474.8987m
R5 2 N5 433.4366m
R6 2 N6 107.3220m
R7 2 N7 1.9771
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820027_2.7n 1 2
C1 1 N7 0.15p
L1 1 N1 2.5n
L2 N1 N2 451.9101p
L3 N2 N3 1.1180n
L4 N3 N4 1.2155n
L5 N4 N5 82.9585p
L6 N5 N6 58.2435p
R1 2 N1 1.1732
R2 2 N2 549.5303m
R3 2 N3 846.4830m
R4 2 N4 743.1445m
R5 2 N5 723.0483m
R6 2 N6 156.6633m
R7 2 N7 1.9708
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820030_3n 1 2
C1 1 N7 0.16p
L1 1 N1 2.7n
L2 N1 N2 444.7303p
L3 N2 N3 1.1012n
L4 N3 N4 1.2155n
L5 N4 N5 83.0034p
L6 N5 N6 58.2841p
R1 2 N1 1.2165
R2 2 N2 436.5621m
R3 2 N3 841.7246m
R4 2 N4 754.1610m
R5 2 N5 734.6394m
R6 2 N6 159.1004m
R7 2 N7 1.9996
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820033_3.3n 1 2
C1 1 N7 0.17p
L1 1 N1 3n
L2 N1 N2 518.9881p
L3 N2 N3 1.1020n
L4 N3 N4 1.2155n
L5 N4 N5 83.0114p
L6 N5 N6 58.2939p
R1 2 N1 1.2395
R2 2 N2 463.4615m
R3 2 N3 842.0645m
R4 2 N4 754.9942m
R5 2 N5 735.5115m
R6 2 N6 159.2744m
R7 2 N7 1.9991
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820036_3.6n 1 2
C1 1 N7 0.17p
L1 1 N1 3.1n
L2 N1 N2 608.2147p
L3 N2 N3 1.1172n
L4 N3 N4 1.2155n
L5 N4 N5 83.1586p
L6 N5 N6 58.4197p
R1 2 N1 1.4984
R2 2 N2 517.4638m
R3 2 N3 854.9344m
R4 2 N4 771.4929m
R5 2 N5 752.4757m
R6 2 N6 162.7767m
R7 2 N7 1.9973
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820039_3.9n 1 2
C1 1 N7 0.18p
L1 1 N1 3.4n
L2 N1 N2 724.0042p
L3 N2 N3 1.2272n
L4 N3 N4 1.2155n
L5 N4 N5 87.5879p
L6 N5 N6 61.4504p
R1 2 N1 1.6668
R2 2 N2 895.5857m
R3 2 N3 1.2222
R4 2 N4 1.0695
R5 2 N5 1.0493
R6 2 N6 224.8339m
R7 2 N7 1.996
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820043_4.3n 1 2
C1 1 N7 0.18p
L1 1 N1 3.8n
L2 N1 N2 536.5024p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 87.6255p
L6 N5 N6 61.4753p
R1 2 N1 1.5631
R2 2 N2 835.3347m
R3 2 N3 1.2226
R4 2 N4 1.0737
R5 2 N5 1.0536
R6 2 N6 225.7728m
R7 2 N7 1.9926
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820047_4.7n 1 2
C1 1 N7 0.19p
L1 1 N1 4.2n
L2 N1 N2 1.0278n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 87.7544p
L6 N5 N6 61.5700p
R1 2 N1 2.0544
R2 2 N2 885.3500m
R3 2 N3 1.2294
R4 2 N4 1.0806
R5 2 N5 1.0604
R6 2 N6 227.1953m
R7 2 N7 1.9893
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820051_5.1n 1 2
C1 1 N7 0.2p
L1 1 N1 4.3n
L2 N1 N2 989.9334p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 87.7832p
L6 N5 N6 61.5911p
R1 2 N1 2.0356
R2 2 N2 872.7899m
R3 2 N3 1.2307
R4 2 N4 1.0824
R5 2 N5 1.0622
R6 2 N6 227.5738m
R7 2 N7 1.9878
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820056_5.6n 1 2
C1 1 N7 0.2p
L1 1 N1 4.8n
L2 N1 N2 810.2328p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 87.9782p
L6 N5 N6 61.7261p
R1 2 N1 1.9768
R2 2 N2 825.7753m
R3 2 N3 1.2417
R4 2 N4 1.0951
R5 2 N5 1.0749
R6 2 N6 230.2620m
R7 2 N7 1.9869
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820062_6.2n 1 2
C1 1 N7 0.23p
L1 1 N1 5.5n
L2 N1 N2 887.9618p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 89.6396p
L6 N5 N6 62.8897p
R1 2 N1 2.2549
R2 2 N2 948.9948m
R3 2 N3 1.3415
R4 2 N4 1.1832
R5 2 N5 1.1619
R6 2 N6 248.6299m
R7 2 N7 1.9848
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820068_6.8n 1 2
C1 1 N7 0.245p
L1 1 N1 6n
L2 N1 N2 986.7214p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 89.7374p
L6 N5 N6 62.9579p
R1 2 N1 2.3076
R2 2 N2 970.8167m
R3 2 N3 1.3472
R4 2 N4 1.1879
R5 2 N5 1.1666
R6 2 N6 249.6103m
R7 2 N7 1.9845
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820075_7.5n 1 2
C1 1 N7 0.26p
L1 1 N1 6.8n
L2 N1 N2 1.1967n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 104.7114p
L6 N5 N6 73.3749p
R1 2 N1 3.1624
R2 2 N2 1.66
R3 2 N3 1.4037
R4 2 N4 1.4122
R5 2 N5 1.4011
R6 2 N6 344.0204m
R7 2 N7 1.9898
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820082_8.2n 1 2
C1 1 N7 0.26p
L1 1 N1 7.3n
L2 N1 N2 1.2338n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 213.2100p
L6 N5 N6 142.1427p
R1 2 N1 3.7067
R2 2 N2 3.7347
R3 2 N3 1.4037
R4 2 N4 1.4122
R5 2 N5 1.4011
R6 2 N6 871.3738m
R7 2 N7 2.4571
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820091_9.1n 1 2
C1 1 N7 0.27p
L1 1 N1 8.5n
L2 N1 N2 1.2338n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 213.2183p
L6 N5 N6 142.1466p
R1 2 N1 3.7067
R2 2 N2 3.7347
R3 2 N3 1.4037
R4 2 N4 1.4122
R5 2 N5 1.4011
R6 2 N6 871.3738m
R7 2 N7 2.4571
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820110_10n 1 2
C1 1 N7 0.3p
L1 1 N1 9n
L2 N1 N2 1.2338n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 213.2276p
L6 N5 N6 142.1511p
R1 2 N1 3.7067
R2 2 N2 3.7347
R3 2 N3 1.4037
R4 2 N4 1.4122
R5 2 N5 1.4011
R6 2 N6 871.3738m
R7 2 N7 2.4572
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820112_12n 1 2
C1 1 N7 0.28p
L1 1 N1 10.5n
L2 N1 N2 1.8094n
L3 N2 N3 2.3114n
L4 N3 N4 2.9882n
L5 N4 N5 223.0101p
L6 N5 N6 146.0117p
R1 2 N1 3.7041
R2 2 N2 3.7312
R3 2 N3 1.4196
R4 2 N4 1.4227
R5 2 N5 1.4107
R6 2 N6 894.6801m
R7 2 N7 19.964
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820115_15n 1 2
C1 1 N7 0.3p
L1 1 N1 13n
L2 N1 N2 2.8900n
L3 N2 N3 2.9360n
L4 N3 N4 4.9211n
L5 N4 N5 233.5643p
L6 N5 N6 150.2062p
R1 2 N1 3.7322
R2 2 N2 3.7245
R3 2 N3 1.445
R4 2 N4 1.4358
R5 2 N5 1.4227
R6 2 N6 922.8717m
R7 2 N7 20.006
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820118_18n 1 2
C1 1 N7 0.3p
L1 1 N1 15n
L2 N1 N2 5.2972n
L3 N2 N3 12.1978n
L4 N3 N4 12.1164n
L5 N4 N5 286.9506p
L6 N5 N6 169.8872p
R1 2 N1 5.2502
R2 2 N2 3.5106
R3 2 N3 1.8337
R4 2 N4 1.4523
R5 2 N5 1.4321
R6 2 N6 938.5966m
R7 2 N7 19.2518
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820122_22n 1 2
C1 1 N7 0.25p
L1 1 N1 18n
L2 N1 N2 4.8135n
L3 N2 N3 12.1901n
L4 N3 N4 12.1164n
L5 N4 N5 313.3623p
L6 N5 N6 179.5176p
R1 2 N1 6.281
R2 2 N2 2.655
R3 2 N3 1.9439
R4 2 N4 1.4591
R5 2 N5 1.4349
R6 2 N6 941.7557m
R7 2 N7 18.6381
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820127_27n 1 2
C1 1 N7 200.9476f
L1 1 N1 26n
L2 N1 N2 8.2024n
L3 N2 N3 104.3551n
L4 N3 N4 119.9382n
L5 N4 N5 340.1304p
L6 N5 N6 211.8392p
R1 2 N1 8.0835
R2 2 N2 2.9012
R3 2 N3 2.1349
R4 2 N4 1.5597
R5 2 N5 1.5371
R6 2 N6 1.1487
R7 2 N7 23.2731
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820133_33n 1 2
C1 1 N7 163.0458f
L1 1 N1 30n
L2 N1 N2 7.1960n
L3 N2 N3 13.7924n
L4 N3 N4 23.4261n
L5 N4 N5 831.4115p
L6 N5 N6 639.4310p
R1 2 N1 12.2013
R2 2 N2 4.2270
R3 2 N3 4.4892
R4 2 N4 4.4448
R5 2 N5 4.4269
R6 2 N6 4.6799
R7 2 N7 29.8567
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840010_1n 1 2
C1 1 N7 303.1247f
L1 1 N1 0.95n
L2 N1 N2 65.2500p
L3 N2 N3 338.7089p
L4 N3 N4 457.9936p
L5 N4 N5 77.2532p
L6 N5 N6 54.4633p
R1 2 N1 328.8877m
R2 2 N2 160.1876m
R3 2 N3 433.2424m
R4 2 N4 392.2436m
R5 2 N5 348.5373m
R6 2 N6 96.5823m
R7 2 N7 1.9658
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840012_1.2n 1 2
C1 1 N7 290.9565f
L1 1 N1 1.1n
L2 N1 N2 60.2748p
L3 N2 N3 325.0993p
L4 N3 N4 453.4185p
L5 N4 N5 77.2258p
L6 N5 N6 54.4464p
R1 2 N1 249.7455m
R2 2 N2 88.2924m
R3 2 N3 427.5731m
R4 2 N4 391.7073m
R5 2 N5 348.2218m
R6 2 N6 96.5632m
R7 2 N7 1.9654
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840015_1.5n 1 2
C1 1 N7 301.5343f
L1 1 N1 1.4n
L2 N1 N2 82.4129p
L3 N2 N3 325.6749p
L4 N3 N4 452.4484p
L5 N4 N5 77.2232p
L6 N5 N6 54.4467p
R1 2 N1 353.8901m
R2 2 N2 171.3700m
R3 2 N3 426.4000m
R4 2 N4 391.8254m
R5 2 N5 348.4714m
R6 2 N6 96.5964m
R7 2 N7 1.9687
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840018_1.8n 1 2
C1 1 N7 398.2805f
L1 1 N1 1.7n
L2 N1 N2 122.5826p
L3 N2 N3 324.8980p
L4 N3 N4 451.9610p
L5 N4 N5 77.2221p
L6 N5 N6 54.4471p
R1 2 N1 401.5882m
R2 2 N2 178.6316m
R3 2 N3 425.6581m
R4 2 N4 391.9128m
R5 2 N5 348.6322m
R6 2 N6 96.6174m
R7 2 N7 1.9707
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840020_2n 1 2
C1 1 N7 0.3518p
L1 1 N1 1.9n
L2 N1 N2 140.7572p
L3 N2 N3 325.0712p
L4 N3 N4 451.9575p
L5 N4 N5 77.2225p
L6 N5 N6 54.4476p
R1 2 N1 411.2266m
R2 2 N2 182.8559m
R3 2 N3 425.6530m
R4 2 N4 391.9293m
R5 2 N5 348.6542m
R6 2 N6 96.6195m
R7 2 N7 1.9709
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840022_2.2n 1 2
C1 1 N7 0.3p
L1 1 N1 2n
L2 N1 N2 194.5174p
L3 N2 N3 337.1053p
L4 N3 N4 456.3147p
L5 N4 N5 77.2551p
L6 N5 N6 54.4693p
R1 2 N1 481.3036m
R2 2 N2 256.1090m
R3 2 N3 429.1584m
R4 2 N4 393.3525m
R5 2 N5 350.1781m
R6 2 N6 96.7944m
R7 2 N7 1.9727
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840027_2.7n 1 2
C1 1 N7 0.25p
L1 1 N1 2.5n
L2 N1 N2 227.5438p
L3 N2 N3 338.0097p
L4 N3 N4 457.0828p
L5 N4 N5 77.2667p
L6 N5 N6 54.4809p
R1 2 N1 482.4065m
R2 2 N2 263.8750m
R3 2 N3 429.1561m
R4 2 N4 393.8922m
R5 2 N5 350.8211m
R6 2 N6 96.8643m
R7 2 N7 1.968
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840030_3n 1 2
C1 1 N7 0.2345p
L1 1 N1 2.7n
L2 N1 N2 216.6071p
L3 N2 N3 453.0084p
L4 N3 N4 539.1771p
L5 N4 N5 77.8524p
L6 N5 N6 54.8452p
R1 2 N1 705.4217m
R2 2 N2 396.4147m
R3 2 N3 471.3275m
R4 2 N4 413.4665m
R5 2 N5 370.0886m
R6 2 N6 99.0340m
R7 2 N7 1.968
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840033_3.3n 1 2
C1 1 N7 0.213p
L1 1 N1 3n
L2 N1 N2 225.4084p
L3 N2 N3 455.4024p
L4 N3 N4 541.7958p
L5 N4 N5 77.8742p
L6 N5 N6 54.8604p
R1 2 N1 697.9905m
R2 2 N2 400.8828m
R3 2 N3 471.7656m
R4 2 N4 414.2939m
R5 2 N5 370.9735m
R6 2 N6 99.1413m
R7 2 N7 1.9669
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840039_3.9n 1 2
C1 1 N7 0.18p
L1 1 N1 3.55n
L2 N1 N2 364.6300p
L3 N2 N3 472.5891p
L4 N3 N4 555.1859p
L5 N4 N5 77.9756p
L6 N5 N6 54.9279p
R1 2 N1 803.2922m
R2 2 N2 424.2183m
R3 2 N3 477.6879m
R4 2 N4 417.6725m
R5 2 N5 374.3669m
R6 2 N6 99.5435m
R7 2 N7 1.9654
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840047_4.7n 1 2
C1 1 N7 0.149p
L1 1 N1 4.35n
L2 N1 N2 473.8107p
L3 N2 N3 530.5532p
L4 N3 N4 600.1689p
L5 N4 N5 78.3015p
L6 N5 N6 55.1354p
R1 2 N1 980.9916m
R2 2 N2 461.4220m
R3 2 N3 499.3521m
R4 2 N4 428.0957m
R5 2 N5 384.5885m
R6 2 N6 100.7801m
R7 2 N7 1.9637
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840056_5.6n 1 2
C1 1 N7 0.16p
L1 1 N1 5.1n
L2 N1 N2 548.0166p
L3 N2 N3 695.2921p
L4 N3 N4 729.9965p
L5 N4 N5 79.2453p
L6 N5 N6 55.7427p
R1 2 N1 1.1969
R2 2 N2 537.6646m
R3 2 N3 560.9455m
R4 2 N4 457.3494m
R5 2 N5 413.1605m
R6 2 N6 104.4004m
R7 2 N7 1.9622
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840068_6.8n 1 2
C1 1 N7 0.2p
L1 1 N1 6.3n
L2 N1 N2 641.3845p
L3 N2 N3 858.6523p
L4 N3 N4 858.3655p
L5 N4 N5 80.1792p
L6 N5 N6 56.3465p
R1 2 N1 1.3589
R2 2 N2 624.6770m
R3 2 N3 619.7612m
R4 2 N4 485.6288m
R5 2 N5 440.8128m
R6 2 N6 108.1890m
R7 2 N7 1.96
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840075_7.5n 1 2
C1 1 N7 0.2p
L1 1 N1 6.9n
L2 N1 N2 774.1596p
L3 N2 N3 973.9145p
L4 N3 N4 958.2757p
L5 N4 N5 80.9143p
L6 N5 N6 56.8263p
R1 2 N1 1.6231
R2 2 N2 662.6402m
R3 2 N3 659.3265m
R4 2 N4 508.1561m
R5 2 N5 463.1075m
R6 2 N6 111.4535m
R7 2 N7 1.9594
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840082_8.2n 1 2
C1 1 N7 0.238p
L1 1 N1 7.5n
L2 N1 N2 872.6976p
L3 N2 N3 1.3379n
L4 N3 N4 1.2702n
L5 N4 N5 83.2046p
L6 N5 N6 58.3299p
R1 2 N1 2.0355
R2 2 N2 774.7286m
R3 2 N3 784.9732m
R4 2 N4 573.8908m
R5 2 N5 527.4021m
R6 2 N6 121.4802m
R7 2 N7 1.9647
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840110_10n 1 2
C1 1 N7 0.247p
L1 1 N1 9n
L2 N1 N2 919.9560p
L3 N2 N3 1.7519n
L4 N3 N4 1.6458n
L5 N4 N5 86.0149p
L6 N5 N6 60.2134p
R1 2 N1 2.4703
R2 2 N2 986.4197m
R3 2 N3 901.7846m
R4 2 N4 654.0942m
R5 2 N5 606.7364m
R6 2 N6 135.1699m
R7 2 N7 1.9965
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840112_12n 1 2
C1 1 N7 200f
L1 1 N1 11n
L2 N1 N2 1.1939n
L3 N2 N3 2.6748n
L4 N3 N4 3.6577n
L5 N4 N5 88.3436p
L6 N5 N6 61.8040p
R1 2 N1 3.1352
R2 2 N2 1.0748
R3 2 N3 988.1124m
R4 2 N4 716.1332m
R5 2 N5 667.4508m
R6 2 N6 224.5649m
R7 2 N7 2.0522
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840115_15n 1 2
C1 1 N7 160.7748f
L1 1 N1 13.5n
L2 N1 N2 1.7873n
L3 N2 N3 4.8391n
L4 N3 N4 4.7907n
L5 N4 N5 88.6137p
L6 N5 N6 62.1276p
R1 2 N1 3.6822
R2 2 N2 1.1151
R3 2 N3 1.0085
R4 2 N4 719.8343m
R5 2 N5 671.0381m
R6 2 N6 238.5628m
R7 2 N7 2.0775
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840118_18n 1 2
C1 1 N7 217.9024f
L1 1 N1 15n
L2 N1 N2 1.9753n
L3 N2 N3 4.8275n
L4 N3 N4 4.7925n
L5 N4 N5 88.6142p
L6 N5 N6 62.1281p
R1 2 N1 3.6961
R2 2 N2 1.1201
R3 2 N3 1.0077
R4 2 N4 719.8707m
R5 2 N5 671.0790m
R6 2 N6 238.8610m
R7 2 N7 2.0819
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840122_22n 1 2
C1 1 N7 200.3328f
L1 1 N1 21n
L2 N1 N2 3.2375n
L3 N2 N3 6.6239n
L4 N3 N4 10.2408n
L5 N4 N5 89.1832p
L6 N5 N6 62.7543p
R1 2 N1 4.0958
R2 2 N2 1.8397
R3 2 N3 1.3426
R4 2 N4 1.2006
R5 2 N5 1.1824
R6 2 N6 1.0241
R7 2 N7 2.9085
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840127_27n 1 2
C1 1 N7 202.1367f
L1 1 N1 26n
L2 N1 N2 5.0909n
L3 N2 N3 7.3272n
L4 N3 N4 11.0453n
L5 N4 N5 89.2233p
L6 N5 N6 62.7680p
R1 2 N1 5.2563
R2 2 N2 1.7971
R3 2 N3 1.4004
R4 2 N4 1.2447
R5 2 N5 1.2276
R6 2 N6 1.0833
R7 2 N7 2.9603
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840133_33n 1 2
C1 1 N7 202.1840f
L1 1 N1 30n
L2 N1 N2 4.8271n
L3 N2 N3 8.6215n
L4 N3 N4 11.6697n
L5 N4 N5 89.2842p
L6 N5 N6 62.8211p
R1 2 N1 5.6036
R2 2 N2 1.8486
R3 2 N3 1.4519
R4 2 N4 1.2754
R5 2 N5 1.2589
R6 2 N6 1.1230
R7 2 N7 2.9934
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840139_39n 1 2
C1 1 N7 198.7636f
L1 1 N1 36.5n
L2 N1 N2 6.4916n
L3 N2 N3 11.1728n
L4 N3 N4 13.1271n
L5 N4 N5 89.3785p
L6 N5 N6 62.8772p
R1 2 N1 6.8429
R2 2 N2 1.9069
R3 2 N3 1.5695
R4 2 N4 1.3392
R5 2 N5 1.3239
R6 2 N6 1.2035
R7 2 N7 3.1542
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840147_47n 1 2
C1 1 N7 162.3308f
L1 1 N1 42n
L2 N1 N2 5.3014n
L3 N2 N3 17.7227n
R1 2 N1 10.0979
R2 2 N2 2.8316
R3 2 N3 1.8068
R7 2 N7 27.1851
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840156_56n 1 2
C1 1 N7 200.6576f
L1 1 N1 50n
L2 N1 N2 7.2081n
L3 N2 N3 21.9340n
R1 2 N1 10.2650
R2 2 N2 3.1395
R3 2 N3 2.3882
R7 2 N7 27.0892
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840168_68n 1 2
C1 1 N7 202.7516f
L1 1 N1 60n
L2 N1 N2 9.0841n
L3 N2 N3 21.9905n
R1 2 N1 10.2847
R2 2 N2 3.1554
R3 2 N3 2.4071
R7 2 N7 27.0775
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840182_82n 1 2
C1 1 N7 276.0361f
L1 1 N1 75n
L2 N1 N2 15.5380n
L3 N2 N3 22.1700n
R1 2 N1 10.3860
R2 2 N2 3.2290
R3 2 N3 2.4324
R7 2 N7 27.0369
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840210_100n 1 2
C1 1 N7 222.4657f
L1 1 N1 90n
L2 N1 N2 15.1215n
L3 N2 N3 48.4709n
R1 2 N1 13.9011
R2 2 N2 3.2684
R3 2 N3 2.4258
R7 2 N7 27.1536
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840212_120n 1 2
C1 1 N7 235.7696f
L1 1 N1 110n
L2 N1 N2 22.4659n
L3 N2 N3 55.4460n
R1 2 N1 15.2303
R2 2 N2 3.2928
R3 2 N3 2.4249
R7 2 N7 27.2334
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840215_150n 1 2
C1 1 N7 311.7086f
L1 1 N1 140n
L2 N1 N2 27.6522n
L3 N2 N3 105.6650n
R1 2 N1 14.4361
R2 2 N2 3.6465
R3 2 N3 2.5250
R7 2 N7 27.7529
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840218_180n 1 2
C1 1 N7 310.6462f
L1 1 N1 160n
L2 N1 N2 36.0640n
L3 N2 N3 150.6717n
R1 2 N1 19.6416
R2 2 N2 4.1564
R3 2 N3 2.7302
R7 2 N7 28.2137
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840222_220n 1 2
C1 1 N7 371.8752f
L1 1 N1 200n
L2 N1 N2 41.1623n
L3 N2 N3 157.3825n
R1 2 N1 18.7886
R2 2 N2 4.2719
R3 2 N3 2.7647
R7 2 N7 28.3247
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840227_270n 1 2
C1 1 N7 484.9586f
L1 1 N1 215n
L2 N1 N2 52.7687n
L3 N2 N3 281.3541n
R1 2 N1 23.6986
R2 2 N2 5.9898
R3 2 N3 3.7695
R7 2 N7 29.4800
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860010_1n 1 2
C1 1 N7 253.3443f
L1 1 N1 0.95n
L2 N1 N2 47.5545p
L3 N2 N3 245.4614p
L4 N3 N4 407.4586p
L5 N4 N5 76.9764p
L6 N5 N6 54.3126p
R1 2 N1 126.8322m
R2 2 N2 54.2116m
R3 2 N3 375.0339m
R4 2 N4 386.4628m
R5 2 N5 345.5001m
R6 2 N6 96.3943m
R7 2 N7 2.0097
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860012_1.2n 1 2
C1 1 N7 0.251p
L1 1 N1 1.15n
L2 N1 N2 52.5510p
L3 N2 N3 241.6526p
L4 N3 N4 404.0145p
L5 N4 N5 76.9589p
L6 N5 N6 54.3074p
R1 2 N1 101.4053m
R2 2 N2 36.3922m
R3 2 N3 373.0195m
R4 2 N4 386.1147m
R5 2 N5 345.3103m
R6 2 N6 96.3736m
R7 2 N7 1.9834
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860015_1.5n 1 2
C1 1 N7 685.7829f
L1 1 N1 1.45n
L2 N1 N2 81.2563p
L3 N2 N3 180.2007p
L4 N3 N4 347.4939p
L5 N4 N5 76.5866p
L6 N5 N6 54.0858p
R1 2 N1 152.2261m
R2 2 N2 42.1481m
R3 2 N3 330.1393m
R4 2 N4 374.8059m
R5 2 N5 335.4430m
R6 2 N6 95.3870m
R7 2 N7 2.0011
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860018_1.8n 1 2
C1 1 N7 591.0353f
L1 1 N1 1.75n
L2 N1 N2 85.1257p
L3 N2 N3 169.7646p
L4 N3 N4 337.7894p
L5 N4 N5 76.5247p
L6 N5 N6 54.0514p
R1 2 N1 198.9241m
R2 2 N2 81.4422m
R3 2 N3 322.9534m
R4 2 N4 373.0357m
R5 2 N5 333.9751m
R6 2 N6 95.2462m
R7 2 N7 1.9912
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860022_2.2n 1 2
C1 1 N7 430.9296f
L1 1 N1 2.1n
L2 N1 N2 90.6138p
L3 N2 N3 171.1093p
L4 N3 N4 337.3436p
L5 N4 N5 76.5364p
L6 N5 N6 54.0647p
R1 2 N1 385.1413m
R2 2 N2 253.7605m
R3 2 N3 320.5267m
R4 2 N4 374.6232m
R5 2 N5 336.1118m
R6 2 N6 95.4982m
R7 2 N7 1.9778
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860027_2.7n 1 2
C1 1 N7 367.3491f
L1 1 N1 2.6n
L2 N1 N2 87.9679p
L3 N2 N3 166.0220p
L4 N3 N4 336.1543p
L5 N4 N5 76.5303p
L6 N5 N6 54.0616p
R1 2 N1 282.7960m
R2 2 N2 229.1314m
R3 2 N3 318.8332m
R4 2 N4 374.5220m
R5 2 N5 336.0884m
R6 2 N6 95.4995m
R7 2 N7 1.9738
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860033_3.3n 1 2
C1 1 N7 378.3170f
L1 1 N1 3.2n
L2 N1 N2 93.0372p
L3 N2 N3 165.7777p
L4 N3 N4 329.7786p
L5 N4 N5 76.5031p
L6 N5 N6 54.0506p
R1 2 N1 467.9102m
R2 2 N2 289.6924m
R3 2 N3 309.3230m
R4 2 N4 374.1067m
R5 2 N5 336.1760m
R6 2 N6 95.5281m
R7 2 N7 1.9743
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860039_3.9n 1 2
C1 1 N7 358.3439f
L1 1 N1 3.8n
L2 N1 N2 96.3316p
L3 N2 N3 210.5324p
L4 N3 N4 329.7447p
L5 N4 N5 76.5145p
L6 N5 N6 54.0656p
R1 2 N1 515.8699m
R2 2 N2 382.8945m
R3 2 N3 312.6760m
R4 2 N4 374.6807m
R5 2 N5 336.9814m
R6 2 N6 95.6116m
R7 2 N7 1.9733
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860047_4.7n 1 2
C1 1 N7 207.4560f
L1 1 N1 4.6n
L2 N1 N2 145.4499p
L3 N2 N3 255.3865p
L4 N3 N4 771.9164p
L5 N4 N5 79.8422p
L6 N5 N6 56.1670p
R1 2 N1 1.3334
R2 2 N2 598.0860m
R3 2 N3 482.1981m
R4 2 N4 517.8190m
R5 2 N5 484.2851m
R6 2 N6 113.2627m
R7 2 N7 1.9646
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860056_5.6n 1 2
C1 1 N7 307.4362f
L1 1 N1 5.5n
L2 N1 N2 150.7699p
L3 N2 N3 347.3696p
L4 N3 N4 775.6217p
L5 N4 N5 79.8818p
L6 N5 N6 56.2038p
R1 2 N1 1.3662
R2 2 N2 701.8177m
R3 2 N3 496.5232m
R4 2 N4 519.9930m
R5 2 N5 486.6436m
R6 2 N6 113.6497m
R7 2 N7 1.9666
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860068_6.8n 1 2
C1 1 N7 203.7456f
L1 1 N1 6.7n
L2 N1 N2 154.3756p
L3 N2 N3 568.0239p
L4 N3 N4 864.0274p
L5 N4 N5 80.5853p
L6 N5 N6 56.6928p
R1 2 N1 1.3864
R2 2 N2 867.1365m
R3 2 N3 541.8865m
R4 2 N4 553.3418m
R5 2 N5 521.0993m
R6 2 N6 119.5569m
R7 2 N7 1.9652
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860082_8.2n 1 2
C1 1 N7 286.7186f
L1 1 N1 8n
L2 N1 N2 383.9763p
L3 N2 N3 577.8613p
L4 N3 N4 877.3471p
L5 N4 N5 80.6939p
L6 N5 N6 56.7711p
R1 2 N1 1.4331
R2 2 N2 885.7530m
R3 2 N3 549.1994m
R4 2 N4 559.0027m
R5 2 N5 526.8871m
R6 2 N6 192.4542m
R7 2 N7 1.9688
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860110_10n 1 2
C1 1 N7 309.1723f
L1 1 N1 9.7n
L2 N1 N2 263.5340p
L3 N2 N3 651.8398p
L4 N3 N4 1.5370n
L5 N4 N5 86.1260p
L6 N5 N6 60.7205p
R1 2 N1 2.661
R2 2 N2 1.4533
R3 2 N3 623.6176m
R4 2 N4 808.4747m
R5 2 N5 779.7481m
R6 2 N6 168.3844m
R7 2 N7 2.1381
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860112_12n 1 2
C1 1 N7 233.5137f
L1 1 N1 11.5n
L2 N1 N2 299.7962p
L3 N2 N3 867.7409p
L4 N3 N4 1.8652n
L5 N4 N5 88.6549p
L6 N5 N6 62.4668p
R1 2 N1 2.902
R2 2 N2 1.5978
R3 2 N3 847.8918m
R4 2 N4 949.0222m
R5 2 N5 921.8727m
R6 2 N6 197.6709m
R7 2 N7 2.213
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860115_15n 1 2
C1 1 N7 281.1867f
L1 1 N1 14.3n
L2 N1 N2 572.0200p
L3 N2 N3 963.8894p
L4 N3 N4 2.7337n
L5 N4 N5 88.7561p
L6 N5 N6 62.5523p
R1 2 N1 3.6582
R2 2 N2 1.2809
R3 2 N3 904.8239m
R4 2 N4 1.0166
R5 2 N5 993.0618m
R6 2 N6 688.9841m
R7 2 N7 2.8354
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860118_18n 1 2
C1 1 N7 257.3203f
L1 1 N1 17.2n
L2 N1 N2 696.3271p
L3 N2 N3 1.3542n
L4 N3 N4 4.5151n
L5 N4 N5 88.8582p
L6 N5 N6 62.6063p
R1 2 N1 3.5568
R2 2 N2 1.718
R3 2 N3 1.0975
R4 2 N4 1.0265
R5 2 N5 1.0028
R6 2 N6 708.5253m
R7 2 N7 2.8376
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860122_22n 1 2
C1 1 N7 271.4170f
L1 1 N1 21n
L2 N1 N2 1.2774n
L3 N2 N3 1.4255n
L4 N3 N4 4.6385n
L5 N4 N5 88.8633p
L6 N5 N6 62.6072p
R1 2 N1 3.6413
R2 2 N2 1.8822
R3 2 N3 1.1205
R4 2 N4 1.0294
R5 2 N5 1.0058
R6 2 N6 714.4343m
R7 2 N7 2.8415
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860127_27n 1 2
C1 1 N7 299.9754f
L1 1 N1 26n
L2 N1 N2 1.7453n
L3 N2 N3 1.5773n
L4 N3 N4 6.2073n
L5 N4 N5 88.9424p
L6 N5 N6 62.6347p
R1 2 N1 3.8221
R2 2 N2 2.0623
R3 2 N3 1.2608
R4 2 N4 1.0535
R5 2 N5 1.0305
R6 2 N6 761.4015m
R7 2 N7 2.9109
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860133_33n 1 2
C1 1 N7 374.2262f
L1 1 N1 32n
L2 N1 N2 1.9679n
L3 N2 N3 1.9125n
L4 N3 N4 8.7532n
L5 N4 N5 88.9295p
L6 N5 N6 62.4757p
R1 2 N1 5.1165
R2 2 N2 2.3014
R3 2 N3 1.6708
R4 2 N4 1.1715
R5 2 N5 1.1523
R6 2 N6 961.9105m
R7 2 N7 3.5954
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860139_39n 1 2
C1 1 N7 260.6304f
L1 1 N1 38n
L2 N1 N2 2.7251n
L3 N2 N3 2.1271n
L4 N3 N4 9.5872n
L5 N4 N5 88.9800p
L6 N5 N6 62.5039p
R1 2 N1 5.1899
R2 2 N2 2.6768
R3 2 N3 1.8217
R4 2 N4 1.1963
R5 2 N5 1.1777
R6 2 N6 997.8156m
R7 2 N7 3.5935
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860147_47n 1 2
C1 1 N7 259.2719f
L1 1 N1 45n
L2 N1 N2 2.9828n
L3 N2 N3 2.9611n
L4 N3 N4 14.9837n
L5 N4 N5 89.2468p
L6 N5 N6 62.5958p
R1 2 N1 7.0459
R2 2 N2 4.1453
R3 2 N3 2.513
R4 2 N4 1.3949
R5 2 N5 1.3801
R6 2 N6 1.2624
R7 2 N7 3.7415
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860156_56n 1 2
C1 1 N7 290.8893f
L1 1 N1 53n
L2 N1 N2 2.4150n
L3 N2 N3 3.9697n
L4 N3 N4 14.3863n
L5 N4 N5 89.2238p
L6 N5 N6 62.5877p
R1 2 N1 10.5389
R2 2 N2 6.13
R3 2 N3 2.7611
R4 2 N4 1.6901
R5 2 N5 1.6813
R6 2 N6 1.6175
R7 2 N7 4.9806
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860168_68n 1 2
C1 1 N7 256.0024f
L1 1 N1 64n
L2 N1 N2 2.9410n
L3 N2 N3 4.6959n
L4 N3 N4 16.3531n
L5 N4 N5 89.3228p
L6 N5 N6 62.6194p
R1 2 N1 10.7465
R2 2 N2 6.8255
R3 2 N3 3.0044
R4 2 N4 1.8345
R5 2 N5 1.8267
R6 2 N6 1.7741
R7 2 N7 4.9791
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860182_82n 1 2
C1 1 N7 324.7846f
L1 1 N1 77n
L2 N1 N2 2.9410n
L3 N2 N3 7.0165n
L4 N3 N4 15.9539n
L5 N4 N5 90.3991p
L6 N5 N6 64.1077p
R1 2 N1 12.9498
R2 2 N2 10.3212
R3 2 N3 2.9058
R4 2 N4 2.309
R5 2 N5 2.3045
R6 2 N6 1.9692
R7 2 N7 5.2736
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860210_100n 1 2
C1 1 N7 271.9311f
L1 1 N1 95n
L2 N1 N2 5.2457n
L3 N2 N3 6.4261n
L4 N3 N4 30.7231n
L5 N4 N5 91.3265p
L6 N5 N6 64.5216p
R1 2 N1 15.2743
R2 2 N2 11.7544
R3 2 N3 4.0939
R4 2 N4 2.5767
R5 2 N5 2.5703
R6 2 N6 1.9921
R7 2 N7 5.5196
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860212_120n 1 2
C1 1 N7 255.9158f
L1 1 N1 110n
L2 N1 N2 7.4140n
L3 N2 N3 6.5099n
L4 N3 N4 33.2158n
L5 N4 N5 91.3461p
L6 N5 N6 64.5474p
R1 2 N1 16.3402
R2 2 N2 12.0112
R3 2 N3 4.0823
R4 2 N4 2.5888
R5 2 N5 2.5825
R6 2 N6 2.0122
R7 2 N7 5.5273
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860215_150n 1 2
C1 1 N7 267.7735f
L1 1 N1 138n
L2 N1 N2 8.2869n
L3 N2 N3 8.6209n
L4 N3 N4 45.8243n
L5 N4 N5 91.3513p
L6 N5 N6 64.5476p
R1 2 N1 20.2757
R2 2 N2 12.0733
R3 2 N3 4.1466
R4 2 N4 2.6159
R5 2 N5 2.6097
R6 2 N6 2.0566
R7 2 N7 5.5623
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860218_180n 1 2
C1 1 N7 326.9390f
L1 1 N1 165n
L2 N1 N2 10.6714n
L3 N2 N3 12.8890n
L4 N3 N4 56.9762n
L5 N4 N5 91.4012p
L6 N5 N6 64.6113p
R1 2 N1 21.3957
R2 2 N2 12.8658
R3 2 N3 4.2535
R4 2 N4 2.6846
R5 2 N5 2.6787
R6 2 N6 2.1653
R7 2 N7 5.5917
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860222_220n 1 2
C1 1 N7 365.3891f
L1 1 N1 195n
L2 N1 N2 14.5252n
L3 N2 N3 19.7771n
L4 N3 N4 91.8753n
L5 N4 N5 91.4051p
L6 N5 N6 64.5974p
R1 2 N1 23.0137
R2 2 N2 13.7886
R3 2 N3 4.4534
R4 2 N4 2.8009
R5 2 N5 2.7955
R6 2 N6 2.3391
R7 2 N7 5.6386
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860227_270n 1 2
C1 1 N7 428.0799f
L1 1 N1 245n
L2 N1 N2 20.5679n
L3 N2 N3 29.6333n
L4 N3 N4 167.1143n
L5 N4 N5 91.4132p
L6 N5 N6 64.5925p
R1 2 N1 23.1403
R2 2 N2 14.3894
R3 2 N3 4.492
R4 2 N4 2.8685
R5 2 N5 2.8633
R6 2 N6 2.4348
R7 2 N7 5.6539
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860233_330n 1 2
C1 1 N7 472.4756f
L1 1 N1 300n
L2 N1 N2 22.0220n
L3 N2 N3 30.1450n
L4 N3 N4 278.3487n
L5 N4 N5 91.4129p
L6 N5 N6 64.5915p
R1 2 N1 23.1572
R2 2 N2 14.8213
R3 2 N3 4.5205
R4 2 N4 2.8632
R5 2 N5 2.8579
R6 2 N6 2.4273
R7 2 N7 5.6537
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860239_390n 1 2
C1 1 N7 455.2490f
L1 1 N1 350n
L2 N1 N2 27.4234n
L3 N2 N3 41.1126n
L4 N3 N4 303.5672n
L5 N4 N5 91.4143p
L6 N5 N6 64.5934p
R1 2 N1 23.1373
R2 2 N2 14.3404
R3 2 N3 4.4915
R4 2 N4 2.8712
R5 2 N5 2.866
R6 2 N6 2.4385
R7 2 N7 5.6544
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860243_430n 1 2
C1 1 N7 501.9212f
L1 1 N1 390n
L2 N1 N2 37.4202n
L3 N2 N3 50.5838n
L4 N3 N4 193.6281n
L5 N4 N5 91.4135p
L6 N5 N6 64.5924p
R1 2 N1 25.5154
R2 2 N2 11.4507
R3 2 N3 4.3738
R4 2 N4 2.9199
R5 2 N5 2.9149
R6 2 N6 2.5059
R7 2 N7 5.6596
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860247_470n 1 2
C1 1 N7 529.6931f
L1 1 N1 420n
L2 N1 N2 45.9830n
L3 N2 N3 60.7206n
L4 N3 N4 351.5059n
L5 N4 N5 91.4232p
L6 N5 N6 64.6054p
R1 2 N1 25.5088
R2 2 N2 11.6916
R3 2 N3 4.3817
R4 2 N4 2.9213
R5 2 N5 2.9163
R6 2 N6 2.5078
R7 2 N7 5.6599
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820010G_1n 1 2
C1 1 N7 252.6464f
L1 1 N1 0.95n
L2 N1 N2 219.3834p
L3 N2 N3 343.0117p
L4 N3 N4 459.3208p
L5 N4 N5 77.2700p
L6 N5 N6 54.4817p
R1 2 N1 453.2257m
R2 2 N2 197.3924m
R3 2 N3 434.9411m
R4 2 N4 392.5233m
R5 2 N5 348.7678m
R6 2 N6 96.5857m
R7 2 N7 1.9655
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820012G_1.2n 1 2
C1 1 N7 0.2p
L1 1 N1 1.15n
L2 N1 N2 247.8759p
L3 N2 N3 343.7710p
L4 N3 N4 460.0589p
L5 N4 N5 77.2770p
L6 N5 N6 54.4873p
R1 2 N1 530.8745m
R2 2 N2 199.8839m
R3 2 N3 435.5468m
R4 2 N4 393.2090m
R5 2 N5 349.5902m
R6 2 N6 96.6861m
R7 2 N7 1.9668
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820015G_1.5n 1 2
C1 1 N7 0.15p
L1 1 N1 1.3n
L2 N1 N2 200.4664p
L3 N2 N3 399.6617p
L4 N3 N4 495.4626p
L5 N4 N5 77.5313p
L6 N5 N6 54.6490p
R1 2 N1 719.2764m
R2 2 N2 344.4866m
R3 2 N3 456.1688m
R4 2 N4 402.5555m
R5 2 N5 359.0284m
R6 2 N6 97.7494m
R7 2 N7 1.9706
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820018G_1.8n 1 2
C1 1 N7 0.14p
L1 1 N1 1.7n
L2 N1 N2 335.7177p
L3 N2 N3 596.4608p
L4 N3 N4 706.6429p
L5 N4 N5 79.1069p
L6 N5 N6 55.6649p
R1 2 N1 825.9598m
R2 2 N2 317.3420m
R3 2 N3 532.8549m
R4 2 N4 460.9317m
R5 2 N5 418.9950m
R6 2 N6 105.2425m
R7 2 N7 1.9764
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820020G_2n 1 2
C1 1 N7 0.16p
L1 1 N1 1.8n
L2 N1 N2 201.6446p
L3 N2 N3 623.6153p
L4 N3 N4 747.7181p
L5 N4 N5 79.4118p
L6 N5 N6 55.8564p
R1 2 N1 593.6751m
R2 2 N2 205.9029m
R3 2 N3 540.5001m
R4 2 N4 473.3010m
R5 2 N5 431.9246m
R6 2 N6 107.1230m
R7 2 N7 1.9727
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820022G_2.2n 1 2
C1 1 N7 0.14p
L1 1 N1 2n
L2 N1 N2 364.2086p
L3 N2 N3 637.5231p
L4 N3 N4 755.6190p
L5 N4 N5 79.4712p
L6 N5 N6 55.8973p
R1 2 N1 742.9116m
R2 2 N2 300.6071m
R3 2 N3 545.9497m
R4 2 N4 474.8793m
R5 2 N5 433.3975m
R6 2 N6 107.3178m
R7 2 N7 1.9758
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820024G_2.4n 1 2
C1 1 N7 0.15p
L1 1 N1 2.2n
L2 N1 N2 379.9885p
L3 N2 N3 637.0462p
L4 N3 N4 755.3142p
L5 N4 N5 79.4707p
L6 N5 N6 55.8982p
R1 2 N1 787.4117m
R2 2 N2 299.8665m
R3 2 N3 545.7213m
R4 2 N4 474.8987m
R5 2 N5 433.4366m
R6 2 N6 107.3220m
R7 2 N7 1.9771
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820027G_2.7n 1 2
C1 1 N7 0.15p
L1 1 N1 2.5n
L2 N1 N2 451.9101p
L3 N2 N3 1.1180n
L4 N3 N4 1.2155n
L5 N4 N5 82.9585p
L6 N5 N6 58.2435p
R1 2 N1 1.1732
R2 2 N2 549.5303m
R3 2 N3 846.4830m
R4 2 N4 743.1445m
R5 2 N5 723.0483m
R6 2 N6 156.6633m
R7 2 N7 1.9708
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820030G_3n 1 2
C1 1 N7 0.16p
L1 1 N1 2.7n
L2 N1 N2 444.7303p
L3 N2 N3 1.1012n
L4 N3 N4 1.2155n
L5 N4 N5 83.0034p
L6 N5 N6 58.2841p
R1 2 N1 1.2165
R2 2 N2 436.5621m
R3 2 N3 841.7246m
R4 2 N4 754.1610m
R5 2 N5 734.6394m
R6 2 N6 159.1004m
R7 2 N7 1.9996
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820033G_3.3n 1 2
C1 1 N7 0.17p
L1 1 N1 3n
L2 N1 N2 518.9881p
L3 N2 N3 1.1020n
L4 N3 N4 1.2155n
L5 N4 N5 83.0114p
L6 N5 N6 58.2939p
R1 2 N1 1.2395
R2 2 N2 463.4615m
R3 2 N3 842.0645m
R4 2 N4 754.9942m
R5 2 N5 735.5115m
R6 2 N6 159.2744m
R7 2 N7 1.9991
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820036G_3.6n 1 2
C1 1 N7 0.17p
L1 1 N1 3.1n
L2 N1 N2 608.2147p
L3 N2 N3 1.1172n
L4 N3 N4 1.2155n
L5 N4 N5 83.1586p
L6 N5 N6 58.4197p
R1 2 N1 1.4984
R2 2 N2 517.4638m
R3 2 N3 854.9344m
R4 2 N4 771.4929m
R5 2 N5 752.4757m
R6 2 N6 162.7767m
R7 2 N7 1.9973
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820039G_3.9n 1 2
C1 1 N7 0.18p
L1 1 N1 3.4n
L2 N1 N2 724.0042p
L3 N2 N3 1.2272n
L4 N3 N4 1.2155n
L5 N4 N5 87.5879p
L6 N5 N6 61.4504p
R1 2 N1 1.6668
R2 2 N2 895.5857m
R3 2 N3 1.2222
R4 2 N4 1.0695
R5 2 N5 1.0493
R6 2 N6 224.8339m
R7 2 N7 1.996
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820043G_4.3n 1 2
C1 1 N7 0.18p
L1 1 N1 3.8n
L2 N1 N2 536.5024p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 87.6255p
L6 N5 N6 61.4753p
R1 2 N1 1.5631
R2 2 N2 835.3347m
R3 2 N3 1.2226
R4 2 N4 1.0737
R5 2 N5 1.0536
R6 2 N6 225.7728m
R7 2 N7 1.9926
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820047G_4.7n 1 2
C1 1 N7 0.19p
L1 1 N1 4.2n
L2 N1 N2 1.0278n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 87.7544p
L6 N5 N6 61.5700p
R1 2 N1 2.0544
R2 2 N2 885.3500m
R3 2 N3 1.2294
R4 2 N4 1.0806
R5 2 N5 1.0604
R6 2 N6 227.1953m
R7 2 N7 1.9893
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820051G_5.1n 1 2
C1 1 N7 0.2p
L1 1 N1 4.3n
L2 N1 N2 989.9334p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 87.7832p
L6 N5 N6 61.5911p
R1 2 N1 2.0356
R2 2 N2 872.7899m
R3 2 N3 1.2307
R4 2 N4 1.0824
R5 2 N5 1.0622
R6 2 N6 227.5738m
R7 2 N7 1.9878
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820056G_5.6n 1 2
C1 1 N7 0.2p
L1 1 N1 4.8n
L2 N1 N2 810.2328p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 87.9782p
L6 N5 N6 61.7261p
R1 2 N1 1.9768
R2 2 N2 825.7753m
R3 2 N3 1.2417
R4 2 N4 1.0951
R5 2 N5 1.0749
R6 2 N6 230.2620m
R7 2 N7 1.9869
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820062G_6.2n 1 2
C1 1 N7 0.23p
L1 1 N1 5.5n
L2 N1 N2 887.9618p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 89.6396p
L6 N5 N6 62.8897p
R1 2 N1 2.2549
R2 2 N2 948.9948m
R3 2 N3 1.3415
R4 2 N4 1.1832
R5 2 N5 1.1619
R6 2 N6 248.6299m
R7 2 N7 1.9848
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820068G_6.8n 1 2
C1 1 N7 0.245p
L1 1 N1 6n
L2 N1 N2 986.7214p
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 89.7374p
L6 N5 N6 62.9579p
R1 2 N1 2.3076
R2 2 N2 970.8167m
R3 2 N3 1.3472
R4 2 N4 1.1879
R5 2 N5 1.1666
R6 2 N6 249.6103m
R7 2 N7 1.9845
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820075G_7.5n 1 2
C1 1 N7 0.26p
L1 1 N1 6.8n
L2 N1 N2 1.1967n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 104.7114p
L6 N5 N6 73.3749p
R1 2 N1 3.1624
R2 2 N2 1.66
R3 2 N3 1.4037
R4 2 N4 1.4122
R5 2 N5 1.4011
R6 2 N6 344.0204m
R7 2 N7 1.9898
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820082G_8.2n 1 2
C1 1 N7 0.26p
L1 1 N1 7.3n
L2 N1 N2 1.2338n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 213.2100p
L6 N5 N6 142.1427p
R1 2 N1 3.7067
R2 2 N2 3.7347
R3 2 N3 1.4037
R4 2 N4 1.4122
R5 2 N5 1.4011
R6 2 N6 871.3738m
R7 2 N7 2.4571
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820091G_9.1n 1 2
C1 1 N7 0.27p
L1 1 N1 8.5n
L2 N1 N2 1.2338n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 213.2183p
L6 N5 N6 142.1466p
R1 2 N1 3.7067
R2 2 N2 3.7347
R3 2 N3 1.4037
R4 2 N4 1.4122
R5 2 N5 1.4011
R6 2 N6 871.3738m
R7 2 N7 2.4571
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820110G_10n 1 2
C1 1 N7 0.3p
L1 1 N1 9n
L2 N1 N2 1.2338n
L3 N2 N3 1.2244n
L4 N3 N4 1.2155n
L5 N4 N5 213.2276p
L6 N5 N6 142.1511p
R1 2 N1 3.7067
R2 2 N2 3.7347
R3 2 N3 1.4037
R4 2 N4 1.4122
R5 2 N5 1.4011
R6 2 N6 871.3738m
R7 2 N7 2.4572
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820112G_12n 1 2
C1 1 N7 0.28p
L1 1 N1 10.5n
L2 N1 N2 1.8094n
L3 N2 N3 2.3114n
L4 N3 N4 2.9882n
L5 N4 N5 223.0101p
L6 N5 N6 146.0117p
R1 2 N1 3.7041
R2 2 N2 3.7312
R3 2 N3 1.4196
R4 2 N4 1.4227
R5 2 N5 1.4107
R6 2 N6 894.6801m
R7 2 N7 19.964
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820115G_15n 1 2
C1 1 N7 0.3p
L1 1 N1 13n
L2 N1 N2 2.8900n
L3 N2 N3 2.9360n
L4 N3 N4 4.9211n
L5 N4 N5 233.5643p
L6 N5 N6 150.2062p
R1 2 N1 3.7322
R2 2 N2 3.7245
R3 2 N3 1.445
R4 2 N4 1.4358
R5 2 N5 1.4227
R6 2 N6 922.8717m
R7 2 N7 20.006
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820118G_18n 1 2
C1 1 N7 0.3p
L1 1 N1 15n
L2 N1 N2 5.2972n
L3 N2 N3 12.1978n
L4 N3 N4 12.1164n
L5 N4 N5 286.9506p
L6 N5 N6 169.8872p
R1 2 N1 5.2502
R2 2 N2 3.5106
R3 2 N3 1.8337
R4 2 N4 1.4523
R5 2 N5 1.4321
R6 2 N6 938.5966m
R7 2 N7 19.2518
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820122G_22n 1 2
C1 1 N7 0.25p
L1 1 N1 18n
L2 N1 N2 4.8135n
L3 N2 N3 12.1901n
L4 N3 N4 12.1164n
L5 N4 N5 313.3623p
L6 N5 N6 179.5176p
R1 2 N1 6.281
R2 2 N2 2.655
R3 2 N3 1.9439
R4 2 N4 1.4591
R5 2 N5 1.4349
R6 2 N6 941.7557m
R7 2 N7 18.6381
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820127G_27n 1 2
C1 1 N7 200.9476f
L1 1 N1 26n
L2 N1 N2 8.2024n
L3 N2 N3 104.3551n
L4 N3 N4 119.9382n
L5 N4 N5 340.1304p
L6 N5 N6 211.8392p
R1 2 N1 8.0835
R2 2 N2 2.9012
R3 2 N3 2.1349
R4 2 N4 1.5597
R5 2 N5 1.5371
R6 2 N6 1.1487
R7 2 N7 23.2731
R8 2 1 10g
.ends 
*******
.subckt 0201_7447820133G_33n 1 2
C1 1 N7 163.0458f
L1 1 N1 30n
L2 N1 N2 7.1960n
L3 N2 N3 13.7924n
L4 N3 N4 23.4261n
L5 N4 N5 831.4115p
L6 N5 N6 639.4310p
R1 2 N1 12.2013
R2 2 N2 4.2270
R3 2 N3 4.4892
R4 2 N4 4.4448
R5 2 N5 4.4269
R6 2 N6 4.6799
R7 2 N7 29.8567
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840010G_1n 1 2
C1 1 N7 303.1247f
L1 1 N1 0.95n
L2 N1 N2 65.2500p
L3 N2 N3 338.7089p
L4 N3 N4 457.9936p
L5 N4 N5 77.2532p
L6 N5 N6 54.4633p
R1 2 N1 328.8877m
R2 2 N2 160.1876m
R3 2 N3 433.2424m
R4 2 N4 392.2436m
R5 2 N5 348.5373m
R6 2 N6 96.5823m
R7 2 N7 1.9658
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840012G_1.2n 1 2
C1 1 N7 290.9565f
L1 1 N1 1.1n
L2 N1 N2 60.2748p
L3 N2 N3 325.0993p
L4 N3 N4 453.4185p
L5 N4 N5 77.2258p
L6 N5 N6 54.4464p
R1 2 N1 249.7455m
R2 2 N2 88.2924m
R3 2 N3 427.5731m
R4 2 N4 391.7073m
R5 2 N5 348.2218m
R6 2 N6 96.5632m
R7 2 N7 1.9654
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840015G_1.5n 1 2
C1 1 N7 301.5343f
L1 1 N1 1.4n
L2 N1 N2 82.4129p
L3 N2 N3 325.6749p
L4 N3 N4 452.4484p
L5 N4 N5 77.2232p
L6 N5 N6 54.4467p
R1 2 N1 353.8901m
R2 2 N2 171.3700m
R3 2 N3 426.4000m
R4 2 N4 391.8254m
R5 2 N5 348.4714m
R6 2 N6 96.5964m
R7 2 N7 1.9687
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840018G_1.8n 1 2
C1 1 N7 398.2805f
L1 1 N1 1.7n
L2 N1 N2 122.5826p
L3 N2 N3 324.8980p
L4 N3 N4 451.9610p
L5 N4 N5 77.2221p
L6 N5 N6 54.4471p
R1 2 N1 401.5882m
R2 2 N2 178.6316m
R3 2 N3 425.6581m
R4 2 N4 391.9128m
R5 2 N5 348.6322m
R6 2 N6 96.6174m
R7 2 N7 1.9707
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840020G_2n 1 2
C1 1 N7 0.3518p
L1 1 N1 1.9n
L2 N1 N2 140.7572p
L3 N2 N3 325.0712p
L4 N3 N4 451.9575p
L5 N4 N5 77.2225p
L6 N5 N6 54.4476p
R1 2 N1 411.2266m
R2 2 N2 182.8559m
R3 2 N3 425.6530m
R4 2 N4 391.9293m
R5 2 N5 348.6542m
R6 2 N6 96.6195m
R7 2 N7 1.9709
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840022G_2.2n 1 2
C1 1 N7 0.3p
L1 1 N1 2n
L2 N1 N2 194.5174p
L3 N2 N3 337.1053p
L4 N3 N4 456.3147p
L5 N4 N5 77.2551p
L6 N5 N6 54.4693p
R1 2 N1 481.3036m
R2 2 N2 256.1090m
R3 2 N3 429.1584m
R4 2 N4 393.3525m
R5 2 N5 350.1781m
R6 2 N6 96.7944m
R7 2 N7 1.9727
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840027G_2.7n 1 2
C1 1 N7 0.25p
L1 1 N1 2.5n
L2 N1 N2 227.5438p
L3 N2 N3 338.0097p
L4 N3 N4 457.0828p
L5 N4 N5 77.2667p
L6 N5 N6 54.4809p
R1 2 N1 482.4065m
R2 2 N2 263.8750m
R3 2 N3 429.1561m
R4 2 N4 393.8922m
R5 2 N5 350.8211m
R6 2 N6 96.8643m
R7 2 N7 1.968
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840030G_3n 1 2
C1 1 N7 0.2345p
L1 1 N1 2.7n
L2 N1 N2 216.6071p
L3 N2 N3 453.0084p
L4 N3 N4 539.1771p
L5 N4 N5 77.8524p
L6 N5 N6 54.8452p
R1 2 N1 705.4217m
R2 2 N2 396.4147m
R3 2 N3 471.3275m
R4 2 N4 413.4665m
R5 2 N5 370.0886m
R6 2 N6 99.0340m
R7 2 N7 1.968
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840033G_3.3n 1 2
C1 1 N7 0.213p
L1 1 N1 3n
L2 N1 N2 225.4084p
L3 N2 N3 455.4024p
L4 N3 N4 541.7958p
L5 N4 N5 77.8742p
L6 N5 N6 54.8604p
R1 2 N1 697.9905m
R2 2 N2 400.8828m
R3 2 N3 471.7656m
R4 2 N4 414.2939m
R5 2 N5 370.9735m
R6 2 N6 99.1413m
R7 2 N7 1.9669
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840039G_3.9n 1 2
C1 1 N7 0.18p
L1 1 N1 3.55n
L2 N1 N2 364.6300p
L3 N2 N3 472.5891p
L4 N3 N4 555.1859p
L5 N4 N5 77.9756p
L6 N5 N6 54.9279p
R1 2 N1 803.2922m
R2 2 N2 424.2183m
R3 2 N3 477.6879m
R4 2 N4 417.6725m
R5 2 N5 374.3669m
R6 2 N6 99.5435m
R7 2 N7 1.9654
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840047G_4.7n 1 2
C1 1 N7 0.149p
L1 1 N1 4.35n
L2 N1 N2 473.8107p
L3 N2 N3 530.5532p
L4 N3 N4 600.1689p
L5 N4 N5 78.3015p
L6 N5 N6 55.1354p
R1 2 N1 980.9916m
R2 2 N2 461.4220m
R3 2 N3 499.3521m
R4 2 N4 428.0957m
R5 2 N5 384.5885m
R6 2 N6 100.7801m
R7 2 N7 1.9637
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840056G_5.6n 1 2
C1 1 N7 0.16p
L1 1 N1 5.1n
L2 N1 N2 548.0166p
L3 N2 N3 695.2921p
L4 N3 N4 729.9965p
L5 N4 N5 79.2453p
L6 N5 N6 55.7427p
R1 2 N1 1.1969
R2 2 N2 537.6646m
R3 2 N3 560.9455m
R4 2 N4 457.3494m
R5 2 N5 413.1605m
R6 2 N6 104.4004m
R7 2 N7 1.9622
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840068G_6.8n 1 2
C1 1 N7 0.2p
L1 1 N1 6.3n
L2 N1 N2 641.3845p
L3 N2 N3 858.6523p
L4 N3 N4 858.3655p
L5 N4 N5 80.1792p
L6 N5 N6 56.3465p
R1 2 N1 1.3589
R2 2 N2 624.6770m
R3 2 N3 619.7612m
R4 2 N4 485.6288m
R5 2 N5 440.8128m
R6 2 N6 108.1890m
R7 2 N7 1.96
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840075G_7.5n 1 2
C1 1 N7 0.2p
L1 1 N1 6.9n
L2 N1 N2 774.1596p
L3 N2 N3 973.9145p
L4 N3 N4 958.2757p
L5 N4 N5 80.9143p
L6 N5 N6 56.8263p
R1 2 N1 1.6231
R2 2 N2 662.6402m
R3 2 N3 659.3265m
R4 2 N4 508.1561m
R5 2 N5 463.1075m
R6 2 N6 111.4535m
R7 2 N7 1.9594
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840082G_8.2n 1 2
C1 1 N7 0.238p
L1 1 N1 7.5n
L2 N1 N2 872.6976p
L3 N2 N3 1.3379n
L4 N3 N4 1.2702n
L5 N4 N5 83.2046p
L6 N5 N6 58.3299p
R1 2 N1 2.0355
R2 2 N2 774.7286m
R3 2 N3 784.9732m
R4 2 N4 573.8908m
R5 2 N5 527.4021m
R6 2 N6 121.4802m
R7 2 N7 1.9647
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840110G_10n 1 2
C1 1 N7 0.247p
L1 1 N1 9n
L2 N1 N2 919.9560p
L3 N2 N3 1.7519n
L4 N3 N4 1.6458n
L5 N4 N5 86.0149p
L6 N5 N6 60.2134p
R1 2 N1 2.4703
R2 2 N2 986.4197m
R3 2 N3 901.7846m
R4 2 N4 654.0942m
R5 2 N5 606.7364m
R6 2 N6 135.1699m
R7 2 N7 1.9965
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840112G_12n 1 2
C1 1 N7 200f
L1 1 N1 11n
L2 N1 N2 1.1939n
L3 N2 N3 2.6748n
L4 N3 N4 3.6577n
L5 N4 N5 88.3436p
L6 N5 N6 61.8040p
R1 2 N1 3.1352
R2 2 N2 1.0748
R3 2 N3 988.1124m
R4 2 N4 716.1332m
R5 2 N5 667.4508m
R6 2 N6 224.5649m
R7 2 N7 2.0522
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840115G_15n 1 2
C1 1 N7 160.7748f
L1 1 N1 13.5n
L2 N1 N2 1.7873n
L3 N2 N3 4.8391n
L4 N3 N4 4.7907n
L5 N4 N5 88.6137p
L6 N5 N6 62.1276p
R1 2 N1 3.6822
R2 2 N2 1.1151
R3 2 N3 1.0085
R4 2 N4 719.8343m
R5 2 N5 671.0381m
R6 2 N6 238.5628m
R7 2 N7 2.0775
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840118G_18n 1 2
C1 1 N7 217.9024f
L1 1 N1 15n
L2 N1 N2 1.9753n
L3 N2 N3 4.8275n
L4 N3 N4 4.7925n
L5 N4 N5 88.6142p
L6 N5 N6 62.1281p
R1 2 N1 3.6961
R2 2 N2 1.1201
R3 2 N3 1.0077
R4 2 N4 719.8707m
R5 2 N5 671.0790m
R6 2 N6 238.8610m
R7 2 N7 2.0819
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840122G_22n 1 2
C1 1 N7 200.3328f
L1 1 N1 21n
L2 N1 N2 3.2375n
L3 N2 N3 6.6239n
L4 N3 N4 10.2408n
L5 N4 N5 89.1832p
L6 N5 N6 62.7543p
R1 2 N1 4.0958
R2 2 N2 1.8397
R3 2 N3 1.3426
R4 2 N4 1.2006
R5 2 N5 1.1824
R6 2 N6 1.0241
R7 2 N7 2.9085
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840127G_27n 1 2
C1 1 N7 202.1367f
L1 1 N1 26n
L2 N1 N2 5.0909n
L3 N2 N3 7.3272n
L4 N3 N4 11.0453n
L5 N4 N5 89.2233p
L6 N5 N6 62.7680p
R1 2 N1 5.2563
R2 2 N2 1.7971
R3 2 N3 1.4004
R4 2 N4 1.2447
R5 2 N5 1.2276
R6 2 N6 1.0833
R7 2 N7 2.9603
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840133G_33n 1 2
C1 1 N7 202.1840f
L1 1 N1 30n
L2 N1 N2 4.8271n
L3 N2 N3 8.6215n
L4 N3 N4 11.6697n
L5 N4 N5 89.2842p
L6 N5 N6 62.8211p
R1 2 N1 5.6036
R2 2 N2 1.8486
R3 2 N3 1.4519
R4 2 N4 1.2754
R5 2 N5 1.2589
R6 2 N6 1.1230
R7 2 N7 2.9934
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840139G_39n 1 2
C1 1 N7 198.7636f
L1 1 N1 36.5n
L2 N1 N2 6.4916n
L3 N2 N3 11.1728n
L4 N3 N4 13.1271n
L5 N4 N5 89.3785p
L6 N5 N6 62.8772p
R1 2 N1 6.8429
R2 2 N2 1.9069
R3 2 N3 1.5695
R4 2 N4 1.3392
R5 2 N5 1.3239
R6 2 N6 1.2035
R7 2 N7 3.1542
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840147G_47n 1 2
C1 1 N7 162.3308f
L1 1 N1 42n
L2 N1 N2 5.3014n
L3 N2 N3 17.7227n
R1 2 N1 10.0979
R2 2 N2 2.8316
R3 2 N3 1.8068
R7 2 N7 27.1851
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840156G_56n 1 2
C1 1 N7 200.6576f
L1 1 N1 50n
L2 N1 N2 7.2081n
L3 N2 N3 21.9340n
R1 2 N1 10.2650
R2 2 N2 3.1395
R3 2 N3 2.3882
R7 2 N7 27.0892
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840168G_68n 1 2
C1 1 N7 202.7516f
L1 1 N1 60n
L2 N1 N2 9.0841n
L3 N2 N3 21.9905n
R1 2 N1 10.2847
R2 2 N2 3.1554
R3 2 N3 2.4071
R7 2 N7 27.0775
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840182G_82n 1 2
C1 1 N7 276.0361f
L1 1 N1 75n
L2 N1 N2 15.5380n
L3 N2 N3 22.1700n
R1 2 N1 10.3860
R2 2 N2 3.2290
R3 2 N3 2.4324
R7 2 N7 27.0369
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840210G_100n 1 2
C1 1 N7 222.4657f
L1 1 N1 90n
L2 N1 N2 15.1215n
L3 N2 N3 48.4709n
R1 2 N1 13.9011
R2 2 N2 3.2684
R3 2 N3 2.4258
R7 2 N7 27.1536
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840212G_120n 1 2
C1 1 N7 235.7696f
L1 1 N1 110n
L2 N1 N2 22.4659n
L3 N2 N3 55.4460n
R1 2 N1 15.2303
R2 2 N2 3.2928
R3 2 N3 2.4249
R7 2 N7 27.2334
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840215G_150n 1 2
C1 1 N7 311.7086f
L1 1 N1 140n
L2 N1 N2 27.6522n
L3 N2 N3 105.6650n
R1 2 N1 14.4361
R2 2 N2 3.6465
R3 2 N3 2.5250
R7 2 N7 27.7529
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840218G_180n 1 2
C1 1 N7 310.6462f
L1 1 N1 160n
L2 N1 N2 36.0640n
L3 N2 N3 150.6717n
R1 2 N1 19.6416
R2 2 N2 4.1564
R3 2 N3 2.7302
R7 2 N7 28.2137
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840222G_220n 1 2
C1 1 N7 371.8752f
L1 1 N1 200n
L2 N1 N2 41.1623n
L3 N2 N3 157.3825n
R1 2 N1 18.7886
R2 2 N2 4.2719
R3 2 N3 2.7647
R7 2 N7 28.3247
R8 2 1 10g
.ends 
*******
.subckt 0402_7447840227G_270n 1 2
C1 1 N7 484.9586f
L1 1 N1 215n
L2 N1 N2 52.7687n
L3 N2 N3 281.3541n
R1 2 N1 23.6986
R2 2 N2 5.9898
R3 2 N3 3.7695
R7 2 N7 29.4800
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860010G_1n 1 2
C1 1 N7 253.3443f
L1 1 N1 0.95n
L2 N1 N2 47.5545p
L3 N2 N3 245.4614p
L4 N3 N4 407.4586p
L5 N4 N5 76.9764p
L6 N5 N6 54.3126p
R1 2 N1 126.8322m
R2 2 N2 54.2116m
R3 2 N3 375.0339m
R4 2 N4 386.4628m
R5 2 N5 345.5001m
R6 2 N6 96.3943m
R7 2 N7 2.0097
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860012G_1.2n 1 2
C1 1 N7 0.251p
L1 1 N1 1.15n
L2 N1 N2 52.5510p
L3 N2 N3 241.6526p
L4 N3 N4 404.0145p
L5 N4 N5 76.9589p
L6 N5 N6 54.3074p
R1 2 N1 101.4053m
R2 2 N2 36.3922m
R3 2 N3 373.0195m
R4 2 N4 386.1147m
R5 2 N5 345.3103m
R6 2 N6 96.3736m
R7 2 N7 1.9834
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860015G_1.5n 1 2
C1 1 N7 685.7829f
L1 1 N1 1.45n
L2 N1 N2 81.2563p
L3 N2 N3 180.2007p
L4 N3 N4 347.4939p
L5 N4 N5 76.5866p
L6 N5 N6 54.0858p
R1 2 N1 152.2261m
R2 2 N2 42.1481m
R3 2 N3 330.1393m
R4 2 N4 374.8059m
R5 2 N5 335.4430m
R6 2 N6 95.3870m
R7 2 N7 2.0011
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860018G_1.8n 1 2
C1 1 N7 591.0353f
L1 1 N1 1.75n
L2 N1 N2 85.1257p
L3 N2 N3 169.7646p
L4 N3 N4 337.7894p
L5 N4 N5 76.5247p
L6 N5 N6 54.0514p
R1 2 N1 198.9241m
R2 2 N2 81.4422m
R3 2 N3 322.9534m
R4 2 N4 373.0357m
R5 2 N5 333.9751m
R6 2 N6 95.2462m
R7 2 N7 1.9912
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860022G_2.2n 1 2
C1 1 N7 430.9296f
L1 1 N1 2.1n
L2 N1 N2 90.6138p
L3 N2 N3 171.1093p
L4 N3 N4 337.3436p
L5 N4 N5 76.5364p
L6 N5 N6 54.0647p
R1 2 N1 385.1413m
R2 2 N2 253.7605m
R3 2 N3 320.5267m
R4 2 N4 374.6232m
R5 2 N5 336.1118m
R6 2 N6 95.4982m
R7 2 N7 1.9778
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860027G_2.7n 1 2
C1 1 N7 367.3491f
L1 1 N1 2.6n
L2 N1 N2 87.9679p
L3 N2 N3 166.0220p
L4 N3 N4 336.1543p
L5 N4 N5 76.5303p
L6 N5 N6 54.0616p
R1 2 N1 282.7960m
R2 2 N2 229.1314m
R3 2 N3 318.8332m
R4 2 N4 374.5220m
R5 2 N5 336.0884m
R6 2 N6 95.4995m
R7 2 N7 1.9738
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860033G_3.3n 1 2
C1 1 N7 378.3170f
L1 1 N1 3.2n
L2 N1 N2 93.0372p
L3 N2 N3 165.7777p
L4 N3 N4 329.7786p
L5 N4 N5 76.5031p
L6 N5 N6 54.0506p
R1 2 N1 467.9102m
R2 2 N2 289.6924m
R3 2 N3 309.3230m
R4 2 N4 374.1067m
R5 2 N5 336.1760m
R6 2 N6 95.5281m
R7 2 N7 1.9743
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860039G_3.9n 1 2
C1 1 N7 358.3439f
L1 1 N1 3.8n
L2 N1 N2 96.3316p
L3 N2 N3 210.5324p
L4 N3 N4 329.7447p
L5 N4 N5 76.5145p
L6 N5 N6 54.0656p
R1 2 N1 515.8699m
R2 2 N2 382.8945m
R3 2 N3 312.6760m
R4 2 N4 374.6807m
R5 2 N5 336.9814m
R6 2 N6 95.6116m
R7 2 N7 1.9733
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860047G_4.7n 1 2
C1 1 N7 207.4560f
L1 1 N1 4.6n
L2 N1 N2 145.4499p
L3 N2 N3 255.3865p
L4 N3 N4 771.9164p
L5 N4 N5 79.8422p
L6 N5 N6 56.1670p
R1 2 N1 1.3334
R2 2 N2 598.0860m
R3 2 N3 482.1981m
R4 2 N4 517.8190m
R5 2 N5 484.2851m
R6 2 N6 113.2627m
R7 2 N7 1.9646
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860056G_5.6n 1 2
C1 1 N7 307.4362f
L1 1 N1 5.5n
L2 N1 N2 150.7699p
L3 N2 N3 347.3696p
L4 N3 N4 775.6217p
L5 N4 N5 79.8818p
L6 N5 N6 56.2038p
R1 2 N1 1.3662
R2 2 N2 701.8177m
R3 2 N3 496.5232m
R4 2 N4 519.9930m
R5 2 N5 486.6436m
R6 2 N6 113.6497m
R7 2 N7 1.9666
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860068G_6.8n 1 2
C1 1 N7 203.7456f
L1 1 N1 6.7n
L2 N1 N2 154.3756p
L3 N2 N3 568.0239p
L4 N3 N4 864.0274p
L5 N4 N5 80.5853p
L6 N5 N6 56.6928p
R1 2 N1 1.3864
R2 2 N2 867.1365m
R3 2 N3 541.8865m
R4 2 N4 553.3418m
R5 2 N5 521.0993m
R6 2 N6 119.5569m
R7 2 N7 1.9652
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860082G_8.2n 1 2
C1 1 N7 286.7186f
L1 1 N1 8n
L2 N1 N2 383.9763p
L3 N2 N3 577.8613p
L4 N3 N4 877.3471p
L5 N4 N5 80.6939p
L6 N5 N6 56.7711p
R1 2 N1 1.4331
R2 2 N2 885.7530m
R3 2 N3 549.1994m
R4 2 N4 559.0027m
R5 2 N5 526.8871m
R6 2 N6 192.4542m
R7 2 N7 1.9688
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860110G_10n 1 2
C1 1 N7 309.1723f
L1 1 N1 9.7n
L2 N1 N2 263.5340p
L3 N2 N3 651.8398p
L4 N3 N4 1.5370n
L5 N4 N5 86.1260p
L6 N5 N6 60.7205p
R1 2 N1 2.661
R2 2 N2 1.4533
R3 2 N3 623.6176m
R4 2 N4 808.4747m
R5 2 N5 779.7481m
R6 2 N6 168.3844m
R7 2 N7 2.1381
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860112G_12n 1 2
C1 1 N7 233.5137f
L1 1 N1 11.5n
L2 N1 N2 299.7962p
L3 N2 N3 867.7409p
L4 N3 N4 1.8652n
L5 N4 N5 88.6549p
L6 N5 N6 62.4668p
R1 2 N1 2.902
R2 2 N2 1.5978
R3 2 N3 847.8918m
R4 2 N4 949.0222m
R5 2 N5 921.8727m
R6 2 N6 197.6709m
R7 2 N7 2.213
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860115G_15n 1 2
C1 1 N7 281.1867f
L1 1 N1 14.3n
L2 N1 N2 572.0200p
L3 N2 N3 963.8894p
L4 N3 N4 2.7337n
L5 N4 N5 88.7561p
L6 N5 N6 62.5523p
R1 2 N1 3.6582
R2 2 N2 1.2809
R3 2 N3 904.8239m
R4 2 N4 1.0166
R5 2 N5 993.0618m
R6 2 N6 688.9841m
R7 2 N7 2.8354
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860118G_18n 1 2
C1 1 N7 257.3203f
L1 1 N1 17.2n
L2 N1 N2 696.3271p
L3 N2 N3 1.3542n
L4 N3 N4 4.5151n
L5 N4 N5 88.8582p
L6 N5 N6 62.6063p
R1 2 N1 3.5568
R2 2 N2 1.718
R3 2 N3 1.0975
R4 2 N4 1.0265
R5 2 N5 1.0028
R6 2 N6 708.5253m
R7 2 N7 2.8376
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860122G_22n 1 2
C1 1 N7 271.4170f
L1 1 N1 21n
L2 N1 N2 1.2774n
L3 N2 N3 1.4255n
L4 N3 N4 4.6385n
L5 N4 N5 88.8633p
L6 N5 N6 62.6072p
R1 2 N1 3.6413
R2 2 N2 1.8822
R3 2 N3 1.1205
R4 2 N4 1.0294
R5 2 N5 1.0058
R6 2 N6 714.4343m
R7 2 N7 2.8415
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860127G_27n 1 2
C1 1 N7 299.9754f
L1 1 N1 26n
L2 N1 N2 1.7453n
L3 N2 N3 1.5773n
L4 N3 N4 6.2073n
L5 N4 N5 88.9424p
L6 N5 N6 62.6347p
R1 2 N1 3.8221
R2 2 N2 2.0623
R3 2 N3 1.2608
R4 2 N4 1.0535
R5 2 N5 1.0305
R6 2 N6 761.4015m
R7 2 N7 2.9109
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860133G_33n 1 2
C1 1 N7 374.2262f
L1 1 N1 32n
L2 N1 N2 1.9679n
L3 N2 N3 1.9125n
L4 N3 N4 8.7532n
L5 N4 N5 88.9295p
L6 N5 N6 62.4757p
R1 2 N1 5.1165
R2 2 N2 2.3014
R3 2 N3 1.6708
R4 2 N4 1.1715
R5 2 N5 1.1523
R6 2 N6 961.9105m
R7 2 N7 3.5954
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860139G_39n 1 2
C1 1 N7 260.6304f
L1 1 N1 38n
L2 N1 N2 2.7251n
L3 N2 N3 2.1271n
L4 N3 N4 9.5872n
L5 N4 N5 88.9800p
L6 N5 N6 62.5039p
R1 2 N1 5.1899
R2 2 N2 2.6768
R3 2 N3 1.8217
R4 2 N4 1.1963
R5 2 N5 1.1777
R6 2 N6 997.8156m
R7 2 N7 3.5935
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860147G_47n 1 2
C1 1 N7 259.2719f
L1 1 N1 45n
L2 N1 N2 2.9828n
L3 N2 N3 2.9611n
L4 N3 N4 14.9837n
L5 N4 N5 89.2468p
L6 N5 N6 62.5958p
R1 2 N1 7.0459
R2 2 N2 4.1453
R3 2 N3 2.513
R4 2 N4 1.3949
R5 2 N5 1.3801
R6 2 N6 1.2624
R7 2 N7 3.7415
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860156G_56n 1 2
C1 1 N7 290.8893f
L1 1 N1 53n
L2 N1 N2 2.4150n
L3 N2 N3 3.9697n
L4 N3 N4 14.3863n
L5 N4 N5 89.2238p
L6 N5 N6 62.5877p
R1 2 N1 10.5389
R2 2 N2 6.13
R3 2 N3 2.7611
R4 2 N4 1.6901
R5 2 N5 1.6813
R6 2 N6 1.6175
R7 2 N7 4.9806
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860168G_68n 1 2
C1 1 N7 256.0024f
L1 1 N1 64n
L2 N1 N2 2.9410n
L3 N2 N3 4.6959n
L4 N3 N4 16.3531n
L5 N4 N5 89.3228p
L6 N5 N6 62.6194p
R1 2 N1 10.7465
R2 2 N2 6.8255
R3 2 N3 3.0044
R4 2 N4 1.8345
R5 2 N5 1.8267
R6 2 N6 1.7741
R7 2 N7 4.9791
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860182G_82n 1 2
C1 1 N7 324.7846f
L1 1 N1 77n
L2 N1 N2 2.9410n
L3 N2 N3 7.0165n
L4 N3 N4 15.9539n
L5 N4 N5 90.3991p
L6 N5 N6 64.1077p
R1 2 N1 12.9498
R2 2 N2 10.3212
R3 2 N3 2.9058
R4 2 N4 2.309
R5 2 N5 2.3045
R6 2 N6 1.9692
R7 2 N7 5.2736
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860210G_100n 1 2
C1 1 N7 271.9311f
L1 1 N1 95n
L2 N1 N2 5.2457n
L3 N2 N3 6.4261n
L4 N3 N4 30.7231n
L5 N4 N5 91.3265p
L6 N5 N6 64.5216p
R1 2 N1 15.2743
R2 2 N2 11.7544
R3 2 N3 4.0939
R4 2 N4 2.5767
R5 2 N5 2.5703
R6 2 N6 1.9921
R7 2 N7 5.5196
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860212G_120n 1 2
C1 1 N7 255.9158f
L1 1 N1 110n
L2 N1 N2 7.4140n
L3 N2 N3 6.5099n
L4 N3 N4 33.2158n
L5 N4 N5 91.3461p
L6 N5 N6 64.5474p
R1 2 N1 16.3402
R2 2 N2 12.0112
R3 2 N3 4.0823
R4 2 N4 2.5888
R5 2 N5 2.5825
R6 2 N6 2.0122
R7 2 N7 5.5273
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860215G_150n 1 2
C1 1 N7 267.7735f
L1 1 N1 138n
L2 N1 N2 8.2869n
L3 N2 N3 8.6209n
L4 N3 N4 45.8243n
L5 N4 N5 91.3513p
L6 N5 N6 64.5476p
R1 2 N1 20.2757
R2 2 N2 12.0733
R3 2 N3 4.1466
R4 2 N4 2.6159
R5 2 N5 2.6097
R6 2 N6 2.0566
R7 2 N7 5.5623
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860218G_180n 1 2
C1 1 N7 326.9390f
L1 1 N1 165n
L2 N1 N2 10.6714n
L3 N2 N3 12.8890n
L4 N3 N4 56.9762n
L5 N4 N5 91.4012p
L6 N5 N6 64.6113p
R1 2 N1 21.3957
R2 2 N2 12.8658
R3 2 N3 4.2535
R4 2 N4 2.6846
R5 2 N5 2.6787
R6 2 N6 2.1653
R7 2 N7 5.5917
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860222G_220n 1 2
C1 1 N7 365.3891f
L1 1 N1 195n
L2 N1 N2 14.5252n
L3 N2 N3 19.7771n
L4 N3 N4 91.8753n
L5 N4 N5 91.4051p
L6 N5 N6 64.5974p
R1 2 N1 23.0137
R2 2 N2 13.7886
R3 2 N3 4.4534
R4 2 N4 2.8009
R5 2 N5 2.7955
R6 2 N6 2.3391
R7 2 N7 5.6386
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860227G_270n 1 2
C1 1 N7 428.0799f
L1 1 N1 245n
L2 N1 N2 20.5679n
L3 N2 N3 29.6333n
L4 N3 N4 167.1143n
L5 N4 N5 91.4132p
L6 N5 N6 64.5925p
R1 2 N1 23.1403
R2 2 N2 14.3894
R3 2 N3 4.492
R4 2 N4 2.8685
R5 2 N5 2.8633
R6 2 N6 2.4348
R7 2 N7 5.6539
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860233G_330n 1 2
C1 1 N7 472.4756f
L1 1 N1 300n
L2 N1 N2 22.0220n
L3 N2 N3 30.1450n
L4 N3 N4 278.3487n
L5 N4 N5 91.4129p
L6 N5 N6 64.5915p
R1 2 N1 23.1572
R2 2 N2 14.8213
R3 2 N3 4.5205
R4 2 N4 2.8632
R5 2 N5 2.8579
R6 2 N6 2.4273
R7 2 N7 5.6537
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860239G_390n 1 2
C1 1 N7 455.2490f
L1 1 N1 350n
L2 N1 N2 27.4234n
L3 N2 N3 41.1126n
L4 N3 N4 303.5672n
L5 N4 N5 91.4143p
L6 N5 N6 64.5934p
R1 2 N1 23.1373
R2 2 N2 14.3404
R3 2 N3 4.4915
R4 2 N4 2.8712
R5 2 N5 2.866
R6 2 N6 2.4385
R7 2 N7 5.6544
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860243G_430n 1 2
C1 1 N7 501.9212f
L1 1 N1 390n
L2 N1 N2 37.4202n
L3 N2 N3 50.5838n
L4 N3 N4 193.6281n
L5 N4 N5 91.4135p
L6 N5 N6 64.5924p
R1 2 N1 25.5154
R2 2 N2 11.4507
R3 2 N3 4.3738
R4 2 N4 2.9199
R5 2 N5 2.9149
R6 2 N6 2.5059
R7 2 N7 5.6596
R8 2 1 10g
.ends 
*******
.subckt 0603_7447860247G_470n 1 2
C1 1 N7 529.6931f
L1 1 N1 420n
L2 N1 N2 45.9830n
L3 N2 N3 60.7206n
L4 N3 N4 351.5059n
L5 N4 N5 91.4232p
L6 N5 N6 64.6054p
R1 2 N1 25.5088
R2 2 N2 11.6916
R3 2 N3 4.3817
R4 2 N4 2.9213
R5 2 N5 2.9163
R6 2 N6 2.5078
R7 2 N7 5.6599
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880015_1.5n 1 2
C1 1 N7 453.7351f
L1 1 N1 1.45n
L2 N1 N2 97.7510p
L3 N2 N3 272.3120p
L4 N3 N4 346.3155p
L5 N4 N5 76.5715p
L6 N5 N6 54.1027p
R1 2 N1 231.6285m
R2 2 N2 86.9697m
R3 2 N3 358.7388m
R4 2 N4 374.9653m
R5 2 N5 335.4371m
R6 2 N6 95.3388m
R7 2 N7 2.0002
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880027_2.7n 1 2
C1 1 N7 370.5358f
L1 1 N1 2.6n
L2 N1 N2 89.2929p
L3 N2 N3 138.7830p
L4 N3 N4 332.2481p
L5 N4 N5 76.5359p
L6 N5 N6 54.0851p
R1 2 N1 324.4136m
R2 2 N2 192.3667m
R3 2 N3 307.5942m
R4 2 N4 374.7480m
R5 2 N5 336.7382m
R6 2 N6 95.5494m
R7 2 N7 1.9562
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880047_4.7n 1 2
C1 1 N7 380.3262f
L1 1 N1 4.6n
L2 N1 N2 62.9873p
L3 N2 N3 189.8775p
L4 N3 N4 770.4824p
L5 N4 N5 79.8434p
L6 N5 N6 56.1732p
R1 2 N1 1.3252
R2 2 N2 569.6958m
R3 2 N3 291.4611m
R4 2 N4 518.3425m
R5 2 N5 484.9844m
R6 2 N6 124.8340m
R7 2 N7 1.9629
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880056_5.6n 1 2
C1 1 N7 417.8944f
L1 1 N1 5.5n
L2 N1 N2 89.9765p
L3 N2 N3 202.8862p
L4 N3 N4 774.3703p
L5 N4 N5 79.9053p
L6 N5 N6 56.2281p
R1 2 N1 1.3445
R2 2 N2 608.0293m
R3 2 N3 448.4145m
R4 2 N4 522.1708m
R5 2 N5 489.3162m
R6 2 N6 156.7441m
R7 2 N7 1.9687
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880068_6.8n 1 2
C1 1 N7 327.6543f
L1 1 N1 6.7n
L2 N1 N2 147.7032p
L3 N2 N3 451.9061p
L4 N3 N4 882.3440p
L5 N4 N5 80.7630p
L6 N5 N6 56.8268p
R1 2 N1 1.3644
R2 2 N2 754.7182m
R3 2 N3 514.5473m
R4 2 N4 565.3774m
R5 2 N5 533.8102m
R6 2 N6 234.4840m
R7 2 N7 1.9655
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880082_8.2n 1 2
C1 1 N7 364.2628f
L1 1 N1 8n
L2 N1 N2 186.9858p
L3 N2 N3 495.2102p
L4 N3 N4 915.0111p
L5 N4 N5 81.0550p
L6 N5 N6 57.0561p
R1 2 N1 1.3571
R2 2 N2 757.3851m
R3 2 N3 545.0157m
R4 2 N4 582.0982m
R5 2 N5 550.8166m
R6 2 N6 322.8298m
R7 2 N7 1.9685
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880110_10n 1 2
C1 1 N7 413.1977f
L1 1 N1 9.7n
L2 N1 N2 148.8577p
L3 N2 N3 252.0940p
L4 N3 N4 943.1212p
L5 N4 N5 86.2628p
L6 N5 N6 60.9923p
R1 2 N1 2.7142
R2 2 N2 1.2388
R3 2 N3 953.8953m
R4 2 N4 863.5495m
R5 2 N5 838.7785m
R6 2 N6 517.8158m
R7 2 N7 2.5106
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880127_27n 1 2
C1 1 N7 478.7462f
L1 1 N1 26n
L2 N1 N2 1.1309n
L3 N2 N3 355.5674p
L4 N3 N4 5.3564n
L5 N4 N5 91.7711p
L6 N5 N6 66.6542p
R1 2 N1 3.2083
R2 2 N2 1.9025
R3 2 N3 1.8277
R4 2 N4 1.1832
R5 2 N5 1.1651
R6 2 N6 973.3438m
R7 2 N7 933.9716m
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880133_33n 1 2
C1 1 N7 425.4063f
L1 1 N1 32n
L2 N1 N2 1.1549n
L3 N2 N3 1.5729n
L4 N3 N4 6.5099n
L5 N4 N5 88.6738p
L6 N5 N6 62.2288p
R1 2 N1 4.9688
R2 2 N2 2.3633
R3 2 N3 1.5105
R4 2 N4 1.1722
R5 2 N5 1.1538
R6 2 N6 964.7568m
R7 2 N7 948.7178m
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880156_56n 1 2
C1 1 N7 497.1717f
L1 1 N1 53n
L2 N1 N2 1.1946n
L3 N2 N3 2.0970n
L4 N3 N4 5.8004n
L5 N4 N5 87.6235p
L6 N5 N6 60.3993p
R1 2 N1 9.5050
R2 2 N2 6.1114
R3 2 N3 2.5141
R4 2 N4 1.7370
R5 2 N5 1.7293
R6 2 N6 1.6696
R7 2 N7 1.3148
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880210_100n 1 2
C1 1 N7 425.5670f
L1 1 N1 95n
L2 N1 N2 4.0949n
L3 N2 N3 779.9348p
L4 N3 N4 9.0957n
L5 N4 N5 91.2600p
L6 N5 N6 64.4001p
R1 2 N1 15.4367
R2 2 N2 11.8692
R3 2 N3 3.8873
R4 2 N4 2.5208
R5 2 N5 2.5141
R6 2 N6 1.8963
R7 2 N7 1.6156
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880212_120n 1 2
C1 1 N7 525.6170f
L1 1 N1 110n
L2 N1 N2 1.4424n
L3 N2 N3 5.7821n
L4 N3 N4 11.6583n
L5 N4 N5 91.3634p
L6 N5 N6 64.4806p
R1 2 N1 15.4856
R2 2 N2 13.2954
R3 2 N3 3.1134
R4 2 N4 2.4554
R5 2 N5 2.4483
R6 2 N6 2.0122
R7 2 N7 5.5273
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880222_220n 1 2
C1 1 N7 515.1440f
L1 1 N1 195n
L2 N1 N2 4.5550n
L3 N2 N3 10.3580n
L4 N3 N4 25.7766n
L5 N4 N5 91.2709p
L6 N5 N6 64.4361p
R1 2 N1 24.6229
R2 2 N2 18.4921
R3 2 N3 4.0010
R4 2 N4 2.8179
R5 2 N5 2.8126
R6 2 N6 2.3636
R7 2 N7 2.4587
R8 2 1 10g
.ends 
*******
.subckt 0805_7447880247_470n 1 2
C1 1 N7 557.0656f
L1 1 N1 420n
L2 N1 N2 24.7521n
L3 N2 N3 35.1655n
L4 N3 N4 267.7875n
L5 N4 N5 91.4235p
L6 N5 N6 64.6063p
R1 2 N1 24.9116
R2 2 N2 10.2555
R3 2 N3 4.3561
R4 2 N4 2.9216
R5 2 N5 2.9166
R6 2 N6 2.5082
R7 2 N7 5.5787
R8 2 1 10g
.ends 
*******










































