**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  SMT Power Inductor
* Matchcode:              WE-LQS
* Library Type:           LTspice
* Version:                rev22b
* Created/modified by:    Ella
* Date and Time:          2022-11-21
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG	
* All Rights Reserved.	
**************************************************	
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy	
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on	
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.	
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.	
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.	
**************************************************	
.subckt 2010_74404020010_1u  1 2
Rp 1 2 1870
Cp 1 2 1.129p
Rs 1 N3 0.094
L1 N3 2 0.724u
.ends 2010_74404020010_1u 
*******
.subckt 2010_74404020015_1.5u  1 2
Rp 1 2 3137
Cp 1 2 1.093p
Rs 1 N3 0.147
L1 N3 2 1.24u
.ends 2010_74404020015_1.5u 
*******
.subckt 2010_74404020022_2.2u  1 2
Rp 1 2 4597
Cp 1 2 1.191p
Rs 1 N3 0.225
L1 N3 2 1.789u
.ends 2010_74404020022_2.2u 
*******
.subckt 2010_74404020033_3.3u  1 2
Rp 1 2 5074
Cp 1 2 1.396p
Rs 1 N3 0.275
L1 N3 2 3.148u
.ends 2010_74404020033_3.3u 
*******
.subckt 2010_74404020047_4.7u  1 2
Rp 1 2 6490
Cp 1 2 1.338p
Rs 1 N3 0.41
L1 N3 2 4.013u
.ends 2010_74404020047_4.7u 
*******
.subckt 2010_74404020068_6.8u  1 2
Rp 1 2 9099
Cp 1 2 1.346p
Rs 1 N3 0.7
L1 N3 2 6.754u
.ends 2010_74404020068_6.8u 
*******
.subckt 2010_74404020100_10u  1 2
Rp 1 2 10056
Cp 1 2 1.922p
Rs 1 N3 0.86
L1 N3 2 9.062u
.ends 2010_74404020100_10u 
*******
.subckt 2010_744040200016_0.16u  1 2
Rp 1 2 425
Cp 1 2 0.67p
Rs 1 N3 0.025
L1 N3 2 0.13u
.ends 2010_744040200016_0.16u 
*******
.subckt 2010_744040200033_0.33u  1 2
Rp 1 2 735
Cp 1 2 0.747p
Rs 1 N3 0.034
L1 N3 2 0.288u
.ends 2010_744040200033_0.33u 
*******
.subckt 2010_744040200047_0.47u  1 2
Rp 1 2 1157
Cp 1 2 0.86p
Rs 1 N3 0.047
L1 N3 2 0.365u
.ends 2010_744040200047_0.47u 
*******
.subckt 2010_744040200068_0.68u  1 2
Rp 1 2 1521
Cp 1 2 1.254p
Rs 1 N3 0.064
L1 N3 2 0.501u
.ends 2010_744040200068_0.68u 
*******
.subckt 2512_74404024010_1u  1 2
Rp 1 2 1713.01
Cp 1 2 1.39575p
Rs 1 N3 0.037
L1 N3 2 1u
.ends 2512_74404024010_1u 
*******
.subckt 2512_74404024015_1.5u  1 2
Rp 1 2 3350.5
Cp 1 2 1.86699p
Rs 1 N3 0.065
L1 N3 2 1.5u
.ends 2512_74404024015_1.5u 
*******
.subckt 2512_74404024022_2.2u  1 2
Rp 1 2 3570.17
Cp 1 2 2.07261p
Rs 1 N3 0.08
L1 N3 2 2.2u
.ends 2512_74404024022_2.2u 
*******
.subckt 2512_74404024033_3.3u  1 2
Rp 1 2 4634.13
Cp 1 2 2.28033p
Rs 1 N3 0.12
L1 N3 2 3.3u
.ends 2512_74404024033_3.3u 
*******
.subckt 2512_74404024047_4.7u  1 2
Rp 1 2 5885.21
Cp 1 2 2.65815p
Rs 1 N3 0.175
L1 N3 2 4.7u
.ends 2512_74404024047_4.7u 
*******
.subckt 2512_74404024068_6.8u  1 2
Rp 1 2 8632.28
Cp 1 2 2.43206p
Rs 1 N3 0.3
L1 N3 2 6.8u
.ends 2512_74404024068_6.8u 
*******
.subckt 2512_74404024100_10u  1 2
Rp 1 2 11069.7
Cp 1 2 2.1441p
Rs 1 N3 0.435
L1 N3 2 10u
.ends 2512_74404024100_10u 
*******
.subckt 2512_74404024101_100u  1 2
Rp 1 2 61437
Cp 1 2 2.189p
Rs 1 N3 4.5
L1 N3 2 109.209u
.ends 2512_74404024101_100u 
*******
.subckt 2512_74404024150_15u  1 2
Rp 1 2 10571.2
Cp 1 2 2.26517p
Rs 1 N3 0.83
L1 N3 2 15u
.ends 2512_74404024150_15u 
*******
.subckt 2512_74404024180_18u  1 2
Rp 1 2 19398.2
Cp 1 2 2.33705p
Rs 1 N3 0.83
L1 N3 2 18u
.ends 2512_74404024180_18u 
*******
.subckt 2512_74404024220_22u  1 2
Rp 1 2 19406.8
Cp 1 2 2.40497p
Rs 1 N3 0.91
L1 N3 2 22u
.ends 2512_74404024220_22u 
*******
.subckt 2512_74404024330_33u  1 2
Rp 1 2 29697.6
Cp 1 2 2.69705p
Rs 1 N3 1.53
L1 N3 2 33u
.ends 2512_74404024330_33u 
*******
.subckt 2512_74404024470_47u  1 2
Rp 1 2 33051
Cp 1 2 3.141p
Rs 1 N3 1.6
L1 N3 2 47u
.ends 2512_74404024470_47u 
*******
.subckt 2512_74404024680_68u  1 2
Rp 1 2 40102
Cp 1 2 2.234p
Rs 1 N3 2.5
L1 N3 2 78.513u
.ends 2512_74404024680_68u 
*******
.subckt 2512_744040240016_0.16u  1 2
Rp 1 2 622.24
Cp 1 2 0.53p
Rs 1 N3 0.016
L1 N3 2 0.16u
.ends 2512_744040240016_0.16u 
*******
.subckt 2512_744040240047_0.47u  1 2
Rp 1 2 1626.69
Cp 1 2 1.09302p
Rs 1 N3 0.032
L1 N3 2 0.47u
.ends 2512_744040240047_0.47u 
*******
.subckt 2512_744040240068_0.68u  1 2
Rp 1 2 1882.65
Cp 1 2 1.41457p
Rs 1 N3 0.035
L1 N3 2 0.68u
.ends 2512_744040240068_0.68u 
*******
.subckt 3012_74404031010A_1u  1 2
Rp 1 2 1474
Cp 1 2 0.815p
Rs 1 N3 31
L1 N3 2 0.73u
.ends 3012_74404031010A_1u 
*******
.subckt 3012_74404031027A_2.7u  1 2
Rp 1 2 3619
Cp 1 2 0.937p
Rs 1 N3 80
L1 N3 2 1.93u
.ends 3012_74404031027A_2.7u 
*******
.subckt 3012_74404031047A_4.7u  1 2
Rp 1 2 5805
Cp 1 2 1.06p
Rs 1 N3 139
L1 N3 2 3.63u
.ends 3012_74404031047A_4.7u 
*******
.subckt 3012_74404031068A_6.8u  1 2
Rp 1 2 7010
Cp 1 2 1.07p
Rs 1 N3 164
L1 N3 2 4.93u
.ends 3012_74404031068A_6.8u 
*******
.subckt 3012_74404031100A_10u  1 2
Rp 1 2 9086
Cp 1 2 1.02p
Rs 1 N3 254
L1 N3 2 7.21u
.ends 3012_74404031100A_10u 
*******
.subckt 3012_74404031150A_15u  1 2
Rp 1 2 14034
Cp 1 2 1.025p
Rs 1 N3 403
L1 N3 2 11.53u
.ends 3012_74404031150A_15u 
*******
.subckt 3012_74404031220A_22u  1 2
Rp 1 2 17806
Cp 1 2 1.173p
Rs 1 N3 524
L1 N3 2 17.646u
.ends 3012_74404031220A_22u 
*******
.subckt 3012_74404031330A_33u  1 2
Rp 1 2 24140
Cp 1 2 1.193p
Rs 1 N3 802
L1 N3 2 24.273u
.ends 3012_74404031330A_33u 
*******
.subckt 3012_74404031470A_47u  1 2
Rp 1 2 33061
Cp 1 2 1.145p
Rs 1 N3 1253
L1 N3 2 36.713u
.ends 3012_74404031470A_47u 
*******
.subckt 3015_74404032010_1u  1 2
Rp 1 2 1774.56
Cp 1 2 1.71977p
Rs 1 N3 0.033
L1 N3 2 1u
.ends 3015_74404032010_1u 
*******
.subckt 3015_74404032015_1.5u  1 2
Rp 1 2 2249.94
Cp 1 2 1.97604p
Rs 1 N3 0.04
L1 N3 2 1.5u
.ends 3015_74404032015_1.5u 
*******
.subckt 3015_74404032022_2.2u  1 2
Rp 1 2 2742.87
Cp 1 2 2.35098p
Rs 1 N3 0.05
L1 N3 2 2.2u
.ends 3015_74404032022_2.2u 
*******
.subckt 3015_74404032033_3.3u  1 2
Rp 1 2 4117
Cp 1 2 1.80801p
Rs 1 N3 0.07
L1 N3 2 3.3u
.ends 3015_74404032033_3.3u 
*******
.subckt 3015_74404032047_4.7u  1 2
Rp 1 2 4847.4
Cp 1 2 2.494p
Rs 1 N3 0.096
L1 N3 2 4.7u
.ends 3015_74404032047_4.7u 
*******
.subckt 3015_74404032068_6.8u  1 2
Rp 1 2 5528.9
Cp 1 2 2.52187p
Rs 1 N3 0.12
L1 N3 2 6.8u
.ends 3015_74404032068_6.8u 
*******
.subckt 3015_74404032100_10u  1 2
Rp 1 2 9125.7
Cp 1 2 2.75432p
Rs 1 N3 0.23
L1 N3 2 10u
.ends 3015_74404032100_10u 
*******
.subckt 3015_74404032101_100u  1 2
Rp 1 2 47900
Cp 1 2 2.28p
Rs 1 N3 2.28
L1 N3 2 100u
.ends 3015_74404032101_100u 
*******
.subckt 3015_74404032150_15u  1 2
Rp 1 2 10875.6
Cp 1 2 3.29482p
Rs 1 N3 0.3
L1 N3 2 15u
.ends 3015_74404032150_15u 
*******
.subckt 3015_74404032220_22u  1 2
Rp 1 2 14300.5
Cp 1 2 3.18927p
Rs 1 N3 0.45
L1 N3 2 22u
.ends 3015_74404032220_22u 
*******
.subckt 3015_74404032330_33u  1 2
Rp 1 2 17543.5
Cp 1 2 3.426p
Rs 1 N3 0.911
L1 N3 2 33u
.ends 3015_74404032330_33u 
*******
.subckt 3015_74404032470_47u  1 2
Rp 1 2 19210
Cp 1 2 3.74p
Rs 1 N3 1.05
L1 N3 2 47u
.ends 3015_74404032470_47u 
*******
.subckt 3015_74404032680_68u  1 2
Rp 1 2 44386
Cp 1 2 1.697p
Rs 1 N3 1.6
L1 N3 2 60.208u
.ends 3015_74404032680_68u 
*******
.subckt 3015_744040320047_0.47u  1 2
Rp 1 2 528.945
Cp 1 2 0.711707p
Rs 1 N3 0.018
L1 N3 2 0.47u
.ends 3015_744040320047_0.47u 
*******
.subckt 4012_74404041010_1u  1 2
Rp 1 2 1977
Cp 1 2 1.191p
Rs 1 N3 0.041
L1 N3 2 1u
.ends 4012_74404041010_1u 
*******
.subckt 4012_74404041033_3.3u  1 2
Rp 1 2 3703
Cp 1 2 2.286p
Rs 1 N3 0.069
L1 N3 2 3.3u
.ends 4012_74404041033_3.3u 
*******
.subckt 4012_74404041047_4.7u  1 2
Rp 1 2 4166
Cp 1 2 2.554p
Rs 1 N3 0.091
L1 N3 2 4.7u
.ends 4012_74404041047_4.7u 
*******
.subckt 4012_74404041100_10u  1 2
Rp 1 2 7002
Cp 1 2 3.18p
Rs 1 N3 0.168
L1 N3 2 10u
.ends 4012_74404041100_10u 
*******
.subckt 4012_74404041101_100u  1 2
Rp 1 2 36368
Cp 1 2 3.945p
Rs 1 N3 1.697
L1 N3 2 100u
.ends 4012_74404041101_100u 
*******
.subckt 4012_74404041220_22u  1 2
Rp 1 2 14500
Cp 1 2 2.05p
Rs 1 N3 0.169
L1 N3 2 21.55u
.ends 4012_74404041220_22u 
*******
.subckt 4012_74404041330_33u  1 2
Rp 1 2 18689
Cp 1 2 3.615p
Rs 1 N3 0.628
L1 N3 2 33u
.ends 4012_74404041330_33u 
*******
.subckt 4012_74404041470_47u  1 2
Rp 1 2 23474
Cp 1 2 3.611p
Rs 1 N3 0.987
L1 N3 2 47u
.ends 4012_74404041470_47u 
*******
.subckt 4012_74404041680_68u  1 2
Rp 1 2 32845
Cp 1 2 3.542p
Rs 1 N3 1.495
L1 N3 2 68u
.ends 4012_74404041680_68u 
*******
.subckt 4012_744040410047_0.47u  1 2
Rp 1 2 759.195
Cp 1 2 0.767p
Rs 1 N3 0.028
L1 N3 2 0.47u
.ends 4012_744040410047_0.47u 
*******
.subckt 4018_74404042010_1u  1 2
Rp 1 2 2231.85
Cp 1 2 2.054p
Rs 1 N3 0.027
L1 N3 2 1u
.ends 4018_74404042010_1u 
*******
.subckt 4018_74404042015_1.5u  1 2
Rp 1 2 2724.08
Cp 1 2 2.32667p
Rs 1 N3 0.031
L1 N3 2 1.5u
.ends 4018_74404042015_1.5u 
*******
.subckt 4018_74404042022_2.2u  1 2
Rp 1 2 3751.82
Cp 1 2 2.5503p
Rs 1 N3 0.042
L1 N3 2 2.2u
.ends 4018_74404042022_2.2u 
*******
.subckt 4018_74404042033_3.3u  1 2
Rp 1 2 4600.61
Cp 1 2 3.1796p
Rs 1 N3 0.055
L1 N3 2 3.3u
.ends 4018_74404042033_3.3u 
*******
.subckt 4018_74404042047_4.7u  1 2
Rp 1 2 5553.94
Cp 1 2 3.00991p
Rs 1 N3 0.07
L1 N3 2 4.7u
.ends 4018_74404042047_4.7u 
*******
.subckt 4018_74404042068_6.8u  1 2
Rp 1 2 6815.98
Cp 1 2 2.93071p
Rs 1 N3 0.098
L1 N3 2 6.8u
.ends 4018_74404042068_6.8u 
*******
.subckt 4018_74404042100_10u  1 2
Rp 1 2 8882.27
Cp 1 2 3.43363p
Rs 1 N3 0.15
L1 N3 2 10u
.ends 4018_74404042100_10u 
*******
.subckt 4018_74404042101_100u  1 2
Rp 1 2 42439
Cp 1 2 4.929p
Rs 1 N3 1.43
L1 N3 2 100u
.ends 4018_74404042101_100u 
*******
.subckt 4018_74404042150_15u  1 2
Rp 1 2 12553.3
Cp 1 2 3.70057p
Rs 1 N3 0.21
L1 N3 2 15u
.ends 4018_74404042150_15u 
*******
.subckt 4018_74404042151_150u  1 2
Rp 1 2 81592
Cp 1 2 4.448p
Rs 1 N3 2.853
L1 N3 2 150u
.ends 4018_74404042151_150u 
*******
.subckt 4018_74404042220_22u  1 2
Rp 1 2 15110.8
Cp 1 2 4.36802p
Rs 1 N3 0.29
L1 N3 2 22u
.ends 4018_74404042220_22u 
*******
.subckt 4018_74404042221_220u  1 2
Rp 1 2 97779
Cp 1 2 5.191p
Rs 1 N3 3.45
L1 N3 2 220u
.ends 4018_74404042221_220u 
*******
.subckt 4018_74404042330_33u  1 2
Rp 1 2 20252.2
Cp 1 2 4.14329p
Rs 1 N3 0.46
L1 N3 2 33u
.ends 4018_74404042330_33u 
*******
.subckt 4018_74404042331_330u  1 2
Rp 1 2 152400
Cp 1 2 4.22p
Rs 1 N3 5.3
L1 N3 2 330u
.ends 4018_74404042331_330u 
*******
.subckt 4018_74404042470_47u  1 2
Rp 1 2 24253.8
Cp 1 2 4.28253p
Rs 1 N3 0.62
L1 N3 2 47u
.ends 4018_74404042470_47u 
*******
.subckt 4018_74404042680_68u  1 2
Rp 1 2 34370
Cp 1 2 5.152p
Rs 1 N3 0.84
L1 N3 2 68u
.ends 4018_74404042680_68u 
*******
.subckt 4018_744040420033_0.33u  1 2
Rp 1 2 784.914
Cp 1 2 1.044p
Rs 1 N3 0.013
L1 N3 2 0.33u
.ends 4018_744040420033_0.33u 
*******
.subckt 4025_74404043010A_1u  1 2
Rp 1 2 1489
Cp 1 2 1.29p
Rs 1 N3 0.014
L1 N3 2 0.639u
.ends 4025_74404043010A_1u 
*******
.subckt 4025_74404043022A_2.2u  1 2
Rp 1 2 3403
Cp 1 2 1.508p
Rs 1 N3 0.023
L1 N3 2 1.464u
.ends 4025_74404043022A_2.2u 
*******
.subckt 4025_74404043033A_3.3u  1 2
Rp 1 2 4904
Cp 1 2 1.655p
Rs 1 N3 0.033
L1 N3 2 2.463u
.ends 4025_74404043033A_3.3u 
*******
.subckt 4025_74404043047A_4.7u  1 2
Rp 1 2 6075
Cp 1 2 1.764p
Rs 1 N3 0.046
L1 N3 2 3.682u
.ends 4025_74404043047A_4.7u 
*******
.subckt 4025_74404043100A_10u  1 2
Rp 1 2 13323
Cp 1 2 1.948p
Rs 1 N3 0.089
L1 N3 2 7.784u
.ends 4025_74404043100A_10u 
*******
.subckt 4025_74404043101A_100u  1 2
Rp 1 2 86036
Cp 1 2 2.373p
Rs 1 N3 1.043
L1 N3 2 86.223u
.ends 4025_74404043101A_100u 
*******
.subckt 4025_74404043102A_1000u  1 2
Rp 1 2 271033
Cp 1 2 2.62p
Rs 1 N3 10.342
L1 N3 2 1025u
.ends 4025_74404043102A_1000u 
*******
.subckt 4025_74404043150A_15u  1 2
Rp 1 2 15713
Cp 1 2 2.312p
Rs 1 N3 0.132
L1 N3 2 11.785u
.ends 4025_74404043150A_15u 
*******
.subckt 4025_74404043151A_150u  1 2
Rp 1 2 150034
Cp 1 2 1.902p
Rs 1 N3 1.634
L1 N3 2 117.883u
.ends 4025_74404043151A_150u 
*******
.subckt 4025_74404043220A_22u  1 2
Rp 1 2 27880
Cp 1 2 1.917p
Rs 1 N3 0.2
L1 N3 2 19.156u
.ends 4025_74404043220A_22u 
*******
.subckt 4025_74404043221A_220u  1 2
Rp 1 2 164796
Cp 1 2 2.493p
Rs 1 N3 2.43
L1 N3 2 200.311u
.ends 4025_74404043221A_220u 
*******
.subckt 4025_74404043330A_33u  1 2
Rp 1 2 32963
Cp 1 2 2.109p
Rs 1 N3 0.316
L1 N3 2 28.373u
.ends 4025_74404043330A_33u 
*******
.subckt 4025_74404043470A_47u  1 2
Rp 1 2 47624
Cp 1 2 2.327p
Rs 1 N3 0.492
L1 N3 2 39.878u
.ends 4025_74404043470A_47u 
*******
.subckt 4025_74404043471A_470u  1 2
Rp 1 2 992355
Cp 1 2 2.412p
Rs 1 N3 3.55
L1 N3 2 420.135u
.ends 4025_74404043471A_470u 
*******
.subckt 5020_74404052010_1u  1 2
Rp 1 2 746
Cp 1 2 3.539p
Rs 1 N3 0.0198
L1 N3 2 1u
.ends 5020_74404052010_1u 
*******
.subckt 5020_74404052012_1.2u  1 2
Rp 1 2 1151.12
Cp 1 2 3.832p
Rs 1 N3 0.0234
L1 N3 2 1.2u
.ends 5020_74404052012_1.2u 
*******
.subckt 5020_74404052015_1.5u  1 2
Rp 1 2 1375.96
Cp 1 2 4.57p
Rs 1 N3 0.0257
L1 N3 2 1.5u
.ends 5020_74404052015_1.5u 
*******
.subckt 5020_74404052022_2.2u  1 2
Rp 1 2 1789
Cp 1 2 4.818p
Rs 1 N3 0.0316
L1 N3 2 2.2u
.ends 5020_74404052022_2.2u 
*******
.subckt 5020_74404052033_3.3u  1 2
Rp 1 2 2582.1
Cp 1 2 4.266p
Rs 1 N3 0.0422
L1 N3 2 3.3u
.ends 5020_74404052033_3.3u 
*******
.subckt 5020_74404052039_3.9u  1 2
Rp 1 2 2489
Cp 1 2 4.171p
Rs 1 N3 0.0505
L1 N3 2 3.9u
.ends 5020_74404052039_3.9u 
*******
.subckt 5020_74404052047_4.7u  1 2
Rp 1 2 3136
Cp 1 2 4.458p
Rs 1 N3 0.0559
L1 N3 2 4.7u
.ends 5020_74404052047_4.7u 
*******
.subckt 5020_74404052056_5.6u  1 2
Rp 1 2 2983
Cp 1 2 7.833p
Rs 1 N3 0.0675
L1 N3 2 5.6u
.ends 5020_74404052056_5.6u 
*******
.subckt 5020_74404052068_6.8u  1 2
Rp 1 2 3076
Cp 1 2 7.38p
Rs 1 N3 0.0827
L1 N3 2 6.8u
.ends 5020_74404052068_6.8u 
*******
.subckt 5020_74404052075_7.5u  1 2
Rp 1 2 4617
Cp 1 2 4.671p
Rs 1 N3 0.0968
L1 N3 2 7.5u
.ends 5020_74404052075_7.5u 
*******
.subckt 5020_74404052100_10u  1 2
Rp 1 2 5418
Cp 1 2 4.975p
Rs 1 N3 0.109
L1 N3 2 10u
.ends 5020_74404052100_10u 
*******
.subckt 5020_74404052101_100u  1 2
Rp 1 2 16782
Cp 1 2 11.992p
Rs 1 N3 1.09
L1 N3 2 100u
.ends 5020_74404052101_100u 
*******
.subckt 5020_74404052150_15u  1 2
Rp 1 2 14175
Cp 1 2 2.244p
Rs 1 N3 0.162
L1 N3 2 13.122u
.ends 5020_74404052150_15u 
*******
.subckt 5020_74404052220_22u  1 2
Rp 1 2 6538
Cp 1 2 11.651p
Rs 1 N3 0.225
L1 N3 2 22u
.ends 5020_74404052220_22u 
*******
.subckt 5020_74404052330_33u  1 2
Rp 1 2 9497
Cp 1 2 10.466p
Rs 1 N3 0.387
L1 N3 2 33u
.ends 5020_74404052330_33u 
*******
.subckt 5020_74404052470_47u  1 2
Rp 1 2 10730
Cp 1 2 11.891p
Rs 1 N3 0.521
L1 N3 2 47u
.ends 5020_74404052470_47u 
*******
.subckt 5020_74404052560_56u  1 2
Rp 1 2 34622
Cp 1 2 2.286p
Rs 1 N3 0.627
L1 N3 2 52.706u
.ends 5020_74404052560_56u 
*******
.subckt 5020_74404052680_68u  1 2
Rp 1 2 14109
Cp 1 2 11.239p
Rs 1 N3 0.627
L1 N3 2 68u
.ends 5020_74404052680_68u 
*******
.subckt 5020_744040520047_0.47u  1 2
Rp 1 2 470
Cp 1 2 2.344p
Rs 1 N3 0.0139
L1 N3 2 0.47u
.ends 5020_744040520047_0.47u 
*******
.subckt 5040_74404054010_1u  1 2
Rp 1 2 2382.76
Cp 1 2 1.05215p
Rs 1 N3 0.012
L1 N3 2 1u
.ends 5040_74404054010_1u 
*******
.subckt 5040_74404054015_1.5u  1 2
Rp 1 2 2903.89
Cp 1 2 1.29794p
Rs 1 N3 0.015
L1 N3 2 1.5u
.ends 5040_74404054015_1.5u 
*******
.subckt 5040_74404054022_2.2u  1 2
Rp 1 2 3313.2
Cp 1 2 2.72661p
Rs 1 N3 0.019
L1 N3 2 2.2u
.ends 5040_74404054022_2.2u 
*******
.subckt 5040_74404054033_3.3u  1 2
Rp 1 2 4741.48
Cp 1 2 4.03036p
Rs 1 N3 0.024
L1 N3 2 3.3u
.ends 5040_74404054033_3.3u 
*******
.subckt 5040_74404054047_4.7u  1 2
Rp 1 2 6232.7
Cp 1 2 4.21371p
Rs 1 N3 0.03
L1 N3 2 4.7u
.ends 5040_74404054047_4.7u 
*******
.subckt 5040_74404054068_6.8u  1 2
Rp 1 2 8059.64
Cp 1 2 4.06082p
Rs 1 N3 0.043
L1 N3 2 6.8u
.ends 5040_74404054068_6.8u 
*******
.subckt 5040_74404054100_10u  1 2
Rp 1 2 11386.7
Cp 1 2 4.55944p
Rs 1 N3 0.064
L1 N3 2 10u
.ends 5040_74404054100_10u 
*******
.subckt 5040_74404054101_100u  1 2
Rp 1 2 38103.4
Cp 1 2 6.18278p
Rs 1 N3 0.56
L1 N3 2 100u
.ends 5040_74404054101_100u 
*******
.subckt 5040_74404054102_1m  1 2
Rp 1 2 358414
Cp 1 2 6.681p
Rs 1 N3 6
L1 N3 2 1000u
.ends 5040_74404054102_1m 
*******
.subckt 5040_74404054150_15u  1 2
Rp 1 2 53628.8
Cp 1 2 5.34333p
Rs 1 N3 0.086
L1 N3 2 15u
.ends 5040_74404054150_15u 
*******
.subckt 5040_74404054151_150u  1 2
Rp 1 2 92731
Cp 1 2 5.524p
Rs 1 N3 0.81
L1 N3 2 131u
.ends 5040_74404054151_150u 
*******
.subckt 5040_74404054220_22u  1 2
Rp 1 2 15968.1
Cp 1 2 4.86858p
Rs 1 N3 0.129
L1 N3 2 22u
.ends 5040_74404054220_22u 
*******
.subckt 5040_74404054221_220u  1 2
Rp 1 2 415855
Cp 1 2 5.846p
Rs 1 N3 1.4
L1 N3 2 209.734u
.ends 5040_74404054221_220u 
*******
.subckt 5040_74404054222_2200u  1 2
Rp 1 2 245560
Cp 1 2 6.44p
Rs 1 N3 12.9
L1 N3 2 2222u
.ends 5040_74404054222_2200u 
*******
.subckt 5040_74404054330_33u  1 2
Rp 1 2 16620.3
Cp 1 2 4.97761p
Rs 1 N3 0.188
L1 N3 2 33u
.ends 5040_74404054330_33u 
*******
.subckt 5040_74404054331_330u  1 2
Rp 1 2 128306
Cp 1 2 8.913p
Rs 1 N3 2.1
L1 N3 2 296.69u
.ends 5040_74404054331_330u 
*******
.subckt 5040_74404054332_3300u  1 2
Rp 1 2 310242
Cp 1 2 10.411p
Rs 1 N3 21.6
L1 N3 2 2430u
.ends 5040_74404054332_3300u 
*******
.subckt 5040_74404054470_47u  1 2
Rp 1 2 23732.6
Cp 1 2 5.67239p
Rs 1 N3 0.272
L1 N3 2 47u
.ends 5040_74404054470_47u 
*******
.subckt 5040_74404054471_470u  1 2
Rp 1 2 81435
Cp 1 2 9.509p
Rs 1 N3 2.95
L1 N3 2 421.19u
.ends 5040_74404054471_470u 
*******
.subckt 5040_74404054680_68u  1 2
Rp 1 2 29490.5
Cp 1 2 5.27529p
Rs 1 N3 0.4
L1 N3 2 68u
.ends 5040_74404054680_68u 
*******
.subckt 5040_74404054681_680u  1 2
Rp 1 2 132164
Cp 1 2 7.357p
Rs 1 N3 3.98
L1 N3 2 665.85u
.ends 5040_74404054681_680u 
*******
.subckt 6028_74404063010_1u  1 2
Rp 1 2 1805.17
Cp 1 2 2.23209p
Rs 1 N3 0.01
L1 N3 2 1u
.ends 6028_74404063010_1u 
*******
.subckt 6028_74404063012_1.2u  1 2
Rp 1 2 2309
Cp 1 2 2.72p
Rs 1 N3 0.011
L1 N3 2 1.2u
.ends 6028_74404063012_1.2u 
*******
.subckt 6028_74404063015_1.5u  1 2
Rp 1 2 2500.45
Cp 1 2 2.48989p
Rs 1 N3 0.013
L1 N3 2 1.5u
.ends 6028_74404063015_1.5u 
*******
.subckt 6028_74404063022_2.2u  1 2
Rp 1 2 4346.53
Cp 1 2 2.85309p
Rs 1 N3 0.02
L1 N3 2 2.2u
.ends 6028_74404063022_2.2u 
*******
.subckt 6028_74404063033_3.3u  1 2
Rp 1 2 5465.48
Cp 1 2 2.78774p
Rs 1 N3 0.025
L1 N3 2 3.3u
.ends 6028_74404063033_3.3u 
*******
.subckt 6028_74404063047_4.7u  1 2
Rp 1 2 6478.1
Cp 1 2 2.9976p
Rs 1 N3 0.03
L1 N3 2 4.7u
.ends 6028_74404063047_4.7u 
*******
.subckt 6028_74404063068_6.8u  1 2
Rp 1 2 8901.72
Cp 1 2 2.9317p
Rs 1 N3 0.047
L1 N3 2 6.8u
.ends 6028_74404063068_6.8u 
*******
.subckt 6028_74404063082_8.2u  1 2
Rp 1 2 10763.8
Cp 1 2 3.17153p
Rs 1 N3 0.055
L1 N3 2 8.2u
.ends 6028_74404063082_8.2u 
*******
.subckt 6028_74404063100_10u  1 2
Rp 1 2 11728.4
Cp 1 2 3.13597p
Rs 1 N3 0.072
L1 N3 2 10u
.ends 6028_74404063100_10u 
*******
.subckt 6028_74404063101_100u  1 2
Rp 1 2 38894.8
Cp 1 2 3.50768p
Rs 1 N3 0.5
L1 N3 2 100u
.ends 6028_74404063101_100u 
*******
.subckt 6028_74404063102_1m  1 2
Rp 1 2 324834
Cp 1 2 6.145p
Rs 1 N3 6.44
L1 N3 2 1000u
.ends 6028_74404063102_1m 
*******
.subckt 6028_74404063150_15u  1 2
Rp 1 2 52665.5
Cp 1 2 3.77615p
Rs 1 N3 0.125
L1 N3 2 15u
.ends 6028_74404063150_15u 
*******
.subckt 6028_74404063220_22u  1 2
Rp 1 2 16563.4
Cp 1 2 3.40651p
Rs 1 N3 0.14
L1 N3 2 22u
.ends 6028_74404063220_22u 
*******
.subckt 6028_74404063330_33u  1 2
Rp 1 2 21914.7
Cp 1 2 3.56615p
Rs 1 N3 0.185
L1 N3 2 33u
.ends 6028_74404063330_33u 
*******
.subckt 6028_74404063470_47u  1 2
Rp 1 2 26736.1
Cp 1 2 3.33866p
Rs 1 N3 0.315
L1 N3 2 47u
.ends 6028_74404063470_47u 
*******
.subckt 6028_74404063680_68u  1 2
Rp 1 2 35422.8
Cp 1 2 3.3614p
Rs 1 N3 0.36
L1 N3 2 68u
.ends 6028_74404063680_68u 
*******
.subckt 6028_74404063681_680u  1 2
Rp 1 2 372702
Cp 1 2 4.61p
Rs 1 N3 5.526
L1 N3 2 723.317u
.ends 6028_74404063681_680u 
*******
.subckt 6028_744040630082_0.82u  1 2
Rp 1 2 1681
Cp 1 2 2.261p
Rs 1 N3 0.01
L1 N3 2 0.82u
.ends 6028_744040630082_0.82u 
*******
.subckt 6045_74404064010_1u  1 2
Rp 1 2 2181.04
Cp 1 2 1.35454p
Rs 1 N3 0.011
L1 N3 2 1u
.ends 6045_74404064010_1u 
*******
.subckt 6045_74404064012_1.2u  1 2
Rp 1 2 2842.9
Cp 1 2 1.65126p
Rs 1 N3 0.01
L1 N3 2 1.2u
.ends 6045_74404064012_1.2u 
*******
.subckt 6045_74404064015_1.5u  1 2
Rp 1 2 2606.14
Cp 1 2 2.12643p
Rs 1 N3 0.012
L1 N3 2 1.5u
.ends 6045_74404064015_1.5u 
*******
.subckt 6045_74404064018_1.8u  1 2
Rp 1 2 3198.37
Cp 1 2 3.20416p
Rs 1 N3 0.012
L1 N3 2 1.8u
.ends 6045_74404064018_1.8u 
*******
.subckt 6045_74404064022_2.2u  1 2
Rp 1 2 4046.34
Cp 1 2 4.18553p
Rs 1 N3 0.014
L1 N3 2 2.2u
.ends 6045_74404064022_2.2u 
*******
.subckt 6045_74404064033_3.3u  1 2
Rp 1 2 5231.48
Cp 1 2 4.34967p
Rs 1 N3 0.021
L1 N3 2 3.3u
.ends 6045_74404064033_3.3u 
*******
.subckt 6045_74404064047_4.7u  1 2
Rp 1 2 7276.7
Cp 1 2 4.75452p
Rs 1 N3 0.026
L1 N3 2 4.7u
.ends 6045_74404064047_4.7u 
*******
.subckt 6045_74404064068_6.8u  1 2
Rp 1 2 9724.71
Cp 1 2 4.99788p
Rs 1 N3 0.031
L1 N3 2 6.8u
.ends 6045_74404064068_6.8u 
*******
.subckt 6045_74404064082_8.2u  1 2
Rp 1 2 11183.8
Cp 1 2 5.54954p
Rs 1 N3 0.043
L1 N3 2 8.2u
.ends 6045_74404064082_8.2u 
*******
.subckt 6045_74404064100_10u  1 2
Rp 1 2 13456.5
Cp 1 2 6.2179p
Rs 1 N3 0.048
L1 N3 2 10u
.ends 6045_74404064100_10u 
*******
.subckt 6045_74404064101_100u  1 2
Rp 1 2 49672.9
Cp 1 2 6.47495p
Rs 1 N3 0.433
L1 N3 2 100u
.ends 6045_74404064101_100u 
*******
.subckt 6045_74404064102_1m  1 2
Rp 1 2 282994
Cp 1 2 6.864p
Rs 1 N3 4.783
L1 N3 2 1000u
.ends 6045_74404064102_1m 
*******
.subckt 6045_74404064120_12u  1 2
Rp 1 2 58118.1
Cp 1 2 7.30919p
Rs 1 N3 0.058
L1 N3 2 12u
.ends 6045_74404064120_12u 
*******
.subckt 6045_74404064121_120u  1 2
Rp 1 2 67827
Cp 1 2 7.536p
Rs 1 N3 0.52
L1 N3 2 120u
.ends 6045_74404064121_120u 
*******
.subckt 6045_74404064150_15u  1 2
Rp 1 2 13176.9
Cp 1 2 6.00805p
Rs 1 N3 0.068
L1 N3 2 15u
.ends 6045_74404064150_15u 
*******
.subckt 6045_74404064151_150u  1 2
Rp 1 2 88382
Cp 1 2 6.917p
Rs 1 N3 0.57
L1 N3 2 150u
.ends 6045_74404064151_150u 
*******
.subckt 6045_74404064152_1.5m  1 2
Rp 1 2 255651
Cp 1 2 10.652p
Rs 1 N3 6.989
L1 N3 2 1500u
.ends 6045_74404064152_1.5m 
*******
.subckt 6045_74404064180_18u  1 2
Rp 1 2 16269.8
Cp 1 2 6.07323p
Rs 1 N3 0.081
L1 N3 2 18u
.ends 6045_74404064180_18u 
*******
.subckt 6045_74404064220_22u  1 2
Rp 1 2 17209.8
Cp 1 2 6.81029p
Rs 1 N3 0.089
L1 N3 2 22u
.ends 6045_74404064220_22u 
*******
.subckt 6045_74404064221_220u  1 2
Rp 1 2 78077
Cp 1 2 8.148p
Rs 1 N3 0.85
L1 N3 2 220u
.ends 6045_74404064221_220u 
*******
.subckt 6045_74404064330_33u  1 2
Rp 1 2 23136.6
Cp 1 2 5.90959p
Rs 1 N3 0.137
L1 N3 2 33u
.ends 6045_74404064330_33u 
*******
.subckt 6045_74404064331_330u  1 2
Rp 1 2 111725
Cp 1 2 7.221p
Rs 1 N3 1.177
L1 N3 2 330u
.ends 6045_74404064331_330u 
*******
.subckt 6045_74404064470_47u  1 2
Rp 1 2 26236.5
Cp 1 2 6.19435p
Rs 1 N3 0.2
L1 N3 2 47u
.ends 6045_74404064470_47u 
*******
.subckt 6045_74404064560_56u  1 2
Rp 1 2 30526
Cp 1 2 11.367p
Rs 1 N3 0.22
L1 N3 2 45.079u
.ends 6045_74404064560_56u 
*******
.subckt 6045_74404064680_68u  1 2
Rp 1 2 32154.2
Cp 1 2 7.6441p
Rs 1 N3 0.289
L1 N3 2 68u
.ends 6045_74404064680_68u 
*******
.subckt 6045_74404064681_680u  1 2
Rp 1 2 117770
Cp 1 2 7.51p
Rs 1 N3 2.1
L1 N3 2 671.67u
.ends 6045_74404064681_680u 
*******
.subckt 6045_744040640047_0.47u  1 2
Rp 1 2 1691
Cp 1 2 1.091p
Rs 1 N3 0.006
L1 N3 2 0.47u
.ends 6045_744040640047_0.47u 
*******
.subckt 6045_744040640068_0.68u  1 2
Rp 1 2 1552
Cp 1 2 1.595p
Rs 1 N3 0.01
L1 N3 2 0.68u
.ends 6045_744040640068_0.68u 
*******
.subckt 8040_74404084010_1u  1 2
Rp 1 2 2123.1
Cp 1 2 1.84879p
Rs 1 N3 0.008
L1 N3 2 1u
.ends 8040_74404084010_1u 
*******
.subckt 8040_74404084015_1.5u  1 2
Rp 1 2 3109.24
Cp 1 2 2.32329p
Rs 1 N3 0.01
L1 N3 2 1.5u
.ends 8040_74404084015_1.5u 
*******
.subckt 8040_74404084022_2.2u  1 2
Rp 1 2 3754.28
Cp 1 2 4.14319p
Rs 1 N3 0.012
L1 N3 2 2.2u
.ends 8040_74404084022_2.2u 
*******
.subckt 8040_74404084033_3.3u  1 2
Rp 1 2 5938.22
Cp 1 2 5.25972p
Rs 1 N3 0.017
L1 N3 2 3.3u
.ends 8040_74404084033_3.3u 
*******
.subckt 8040_74404084047_4.7u  1 2
Rp 1 2 6853.85
Cp 1 2 5.78901p
Rs 1 N3 0.019
L1 N3 2 4.7u
.ends 8040_74404084047_4.7u 
*******
.subckt 8040_74404084068_6.8u  1 2
Rp 1 2 9486.38
Cp 1 2 5.60607p
Rs 1 N3 0.024
L1 N3 2 6.8u
.ends 8040_74404084068_6.8u 
*******
.subckt 8040_74404084082_8.2u  1 2
Rp 1 2 11620.5
Cp 1 2 5.94956p
Rs 1 N3 0.026
L1 N3 2 8.2u
.ends 8040_74404084082_8.2u 
*******
.subckt 8040_74404084100_10u  1 2
Rp 1 2 11946.9
Cp 1 2 5.37055p
Rs 1 N3 0.029
L1 N3 2 10u
.ends 8040_74404084100_10u 
*******
.subckt 8040_74404084101_100u  1 2
Rp 1 2 46943.9
Cp 1 2 6.3045p
Rs 1 N3 0.29
L1 N3 2 100u
.ends 8040_74404084101_100u 
*******
.subckt 8040_74404084102_1m  1 2
Rp 1 2 233948
Cp 1 2 7.1p
Rs 1 N3 2.87
L1 N3 2 1000u
.ends 8040_74404084102_1m 
*******
.subckt 8040_74404084120_12u  1 2
Rp 1 2 53057.6
Cp 1 2 6.72576p
Rs 1 N3 0.04
L1 N3 2 12u
.ends 8040_74404084120_12u 
*******
.subckt 8040_74404084121_120u  1 2
Rp 1 2 58710
Cp 1 2 6.795p
Rs 1 N3 0.347
L1 N3 2 120u
.ends 8040_74404084121_120u 
*******
.subckt 8040_74404084150_15u  1 2
Rp 1 2 15418.7
Cp 1 2 5.75566p
Rs 1 N3 0.047
L1 N3 2 15u
.ends 8040_74404084150_15u 
*******
.subckt 8040_74404084151_150u  1 2
Rp 1 2 83286
Cp 1 2 7.01p
Rs 1 N3 0.478
L1 N3 2 150u
.ends 8040_74404084151_150u 
*******
.subckt 8040_74404084180_18u  1 2
Rp 1 2 16468.2
Cp 1 2 5.8282p
Rs 1 N3 0.053
L1 N3 2 18u
.ends 8040_74404084180_18u 
*******
.subckt 8040_74404084220_22u  1 2
Rp 1 2 19840.6
Cp 1 2 6.46916p
Rs 1 N3 0.069
L1 N3 2 22u
.ends 8040_74404084220_22u 
*******
.subckt 8040_74404084221_220u  1 2
Rp 1 2 105122
Cp 1 2 6.794p
Rs 1 N3 0.592
L1 N3 2 220u
.ends 8040_74404084221_220u 
*******
.subckt 8040_74404084330_33u  1 2
Rp 1 2 20204.8
Cp 1 2 5.65113p
Rs 1 N3 0.097
L1 N3 2 33u
.ends 8040_74404084330_33u 
*******
.subckt 8040_74404084331_330u  1 2
Rp 1 2 142263
Cp 1 2 6.937p
Rs 1 N3 0.865
L1 N3 2 330u
.ends 8040_74404084331_330u 
*******
.subckt 8040_74404084470_47u  1 2
Rp 1 2 24457.1
Cp 1 2 7.00455p
Rs 1 N3 0.136
L1 N3 2 47u
.ends 8040_74404084470_47u 
*******
.subckt 8040_74404084560_56u 1 2
Rp 1 2 27870
Cp 1 2 7.9p
Rs 1 N3 0.18
L1 N3 2 51.4u
.ends 8040_74404084560_56u
*******
.subckt 8040_74404084680_68u  1 2
Rp 1 2 35638.3
Cp 1 2 6.31246p
Rs 1 N3 0.196
L1 N3 2 68u
.ends 8040_74404084680_68u 
*******
.subckt 8040_74404084681_680u  1 2
Rp 1 2 214913
Cp 1 2 5.919p
Rs 1 N3 2.032
L1 N3 2 723.53u
.ends 8040_74404084681_680u 
*******
.subckt 8065_74404086101_100u  1 2
Rp 1 2 49550
Cp 1 2 15.52p
Rs 1 N3 0.238
L1 N3 2 94.56u
.ends 8065_74404086101_100u 
*******
.subckt 8065_74404086102_1000u  1 2
Rp 1 2 129750
Cp 1 2 13.55p
Rs 1 N3 2.35
L1 N3 2 948u
.ends 8065_74404086102_1000u 
*******
.subckt 8065_74404086103_10000u  1 2
Rp 1 2 443000
Cp 1 2 17.65p
Rs 1 N3 22.8
L1 N3 2 8836u
.ends 8065_74404086103_10000u 
*******
.subckt 8065_74404086151_150u  1 2
Rp 1 2 66107
Cp 1 2 15.97p
Rs 1 N3 0.355
L1 N3 2 139.75u
.ends 8065_74404086151_150u 
*******
.subckt 8065_74404086152_1500u  1 2
Rp 1 2 155000
Cp 1 2 14.95p
Rs 1 N3 3.65
L1 N3 2 1429u
.ends 8065_74404086152_1500u 
*******
.subckt 8065_74404086221_220u  1 2
Rp 1 2 90000
Cp 1 2 15.7p
Rs 1 N3 0.555
L1 N3 2 212u
.ends 8065_74404086221_220u 
*******
.subckt 8065_74404086222_2200u  1 2
Rp 1 2 311380
Cp 1 2 10.87p
Rs 1 N3 5
L1 N3 2 2144u
.ends 8065_74404086222_2200u 
*******
.subckt 8065_74404086331_330u  1 2
Rp 1 2 93840
Cp 1 2 14.79p
Rs 1 N3 0.7
L1 N3 2 310.97u
.ends 8065_74404086331_330u 
*******
.subckt 8065_74404086332_3300u  1 2
Rp 1 2 255000
Cp 1 2 15.024p
Rs 1 N3 7.3
L1 N3 2 3069u
.ends 8065_74404086332_3300u 
*******
.subckt 8065_74404086471_470u  1 2
Rp 1 2 106610
Cp 1 2 16.92p
Rs 1 N3 1.2
L1 N3 2 493.31u
.ends 8065_74404086471_470u 
*******
.subckt 8065_74404086472_4700u  1 2
Rp 1 2 371271
Cp 1 2 14.816p
Rs 1 N3 12.15
L1 N3 2 4430u
.ends 8065_74404086472_4700u 
*******
.subckt 8065_74404086681_680u  1 2
Rp 1 2 109785
Cp 1 2 14.707p
Rs 1 N3 1.65
L1 N3 2 651.45u
.ends 8065_74404086681_680u 
*******
.subckt 8065_74404086682_6800u  1 2
Rp 1 2 791553
Cp 1 2 12.992p
Rs 1 N3 18.7
L1 N3 2 6536u
.ends 8065_74404086682_6800u 
*******
