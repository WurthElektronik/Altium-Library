**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Polymer Capacitors
* Matchcode:             WCAP-PTHR
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 870055673001_10uF 1 2
Rser 1 3 0.0214027298475
Lser 2 4 2.934706957E-09
C1 3 4 0.00001
Rpar 3 4 350000
.ends 870055673001_10uF
*******
.subckt 870055673002_22uF 1 2
Rser 1 3 0.00993446943878
Lser 2 4 3.273498602E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 870055673002_22uF
*******
.subckt 870055674003_33uF 1 2
Rser 1 3 0.0107728199644
Lser 2 4 3.157117958E-09
C1 3 4 0.000033
Rpar 3 4 151515.151515152
.ends 870055674003_33uF
*******
.subckt 870055674004_39uF 1 2
Rser 1 3 0.0103409086413
Lser 2 4 3.185369302E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 870055674004_39uF
*******
.subckt 870055674005_47uF 1 2
Rser 1 3 0.0125699233915
Lser 2 4 4.534908902E-09
C1 3 4 0.000047
Rpar 3 4 106382.978723404
.ends 870055674005_47uF
*******
.subckt 870055674006_56uF 1 2
Rser 1 3 0.0094747493131
Lser 2 4 4.207387253E-09
C1 3 4 0.000056
Rpar 3 4 89285.7142857143
.ends 870055674006_56uF
*******
.subckt 870055674007_68uF 1 2
Rser 1 3 0.0130784816817
Lser 2 4 3.439429115E-09
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 870055674007_68uF
*******
.subckt 870055675008_82uF 1 2
Rser 1 3 0.00944800546273
Lser 2 4 7.050474676E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 870055675008_82uF
*******
.subckt 870055675009_100uF 1 2
Rser 1 3 0.0136476609813
Lser 2 4 9.36146617836E-09
C1 3 4 0.0001
Rpar 3 4 50000
.ends 870055675009_100uF
*******
.subckt 870055675010_150uF 1 2
Rser 1 3 0.0130332413108
Lser 2 4 8.803410584E-09
C1 3 4 0.00015
Rpar 3 4 33333.3333333333
.ends 870055675010_150uF
*******
.subckt 870055774001_10uF 1 2
Rser 1 3 0.014424848722
Lser 2 4 7.209081727E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 870055774001_10uF
*******
.subckt 870055774002_22uF 1 2
Rser 1 3 0.014337014827
Lser 2 4 4.619666181E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 870055774002_22uF
*******
.subckt 870055775003_33uF 1 2
Rser 1 3 0.0105908634443
Lser 2 4 5.226495698E-09
C1 3 4 0.000033
Rpar 3 4 151515.151515152
.ends 870055775003_33uF
*******
.subckt 870055775004_39uF 1 2
Rser 1 3 0.0114530926154
Lser 2 4 6.208486852E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 870055775004_39uF
*******
.subckt 870055775005_47uF 1 2
Rser 1 3 0.0109989724954
Lser 2 4 5.350352123E-09
C1 3 4 0.000047
Rpar 3 4 106382.978723404
.ends 870055775005_47uF
*******
.subckt 870055775006_56uF 1 2
Rser 1 3 0.0108800835115
Lser 2 4 6.692979159E-09
C1 3 4 0.000056
Rpar 3 4 89285.7142857143
.ends 870055775006_56uF
*******
.subckt 870055775007_68uF 1 2
Rser 1 3 0.0142844211564
Lser 2 4 6.123867279E-09
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 870055775007_68uF
*******
.subckt 870055874001_10uF 1 2
Rser 1 3 0.0142844211564
Lser 2 4 6.123867279E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 870055874001_10uF
*******
.subckt 870055874002_22uF 1 2
Rser 1 3 0.0133164248124
Lser 2 4 5.014984862E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 870055874002_22uF
*******
.subckt 870055875003_33uF 1 2
Rser 1 3 0.0150612320095
Lser 2 4 7.978889804E-09
C1 3 4 0.000033
Rpar 3 4 151515.151515152
.ends 870055875003_33uF
*******
.subckt 870055875004_39uF 1 2
Rser 1 3 0.0130724870155
Lser 2 4 7.594165845E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 870055875004_39uF
*******
.subckt 870055875005_47uF 1 2
Rser 1 3 0.0123344782098
Lser 2 4 7.380398682E-09
C1 3 4 0.000047
Rpar 3 4 106382.978723404
.ends 870055875005_47uF
*******
.subckt 870055875006_56uF 1 2
Rser 1 3 0.010355477926
Lser 2 4 7.04716567E-09
C1 3 4 0.000056
Rpar 3 4 89285.7142857143
.ends 870055875006_56uF
*******
.subckt 870055974001_10uF 1 2
Rser 1 3 0.0107913922353
Lser 2 4 4.982623278E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 870055974001_10uF
*******
.subckt 870055975002_22uF 1 2
Rser 1 3 0.0108478478375
Lser 2 4 4.312574498E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 870055975002_22uF
*******
.subckt 870055975003_33uF 1 2
Rser 1 3 0.0143277522691
Lser 2 4 6.416844946E-09
C1 3 4 0.000033
Rpar 3 4 151515.151515152
.ends 870055975003_33uF
*******
.subckt 870055975004_47uF 1 2
Rser 1 3 0.0100454268693
Lser 2 4 5.608800366E-09
C1 3 4 0.000047
Rpar 3 4 106382.978723404
.ends 870055975004_47uF
*******
.subckt 870056174001_10uF 1 2
Rser 1 3 0.0122147969484
Lser 2 4 3.967868679E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 870056174001_10uF
*******
.subckt 870056174002_12uF 1 2
Rser 1 3 0.0127666247444
Lser 2 4 6.575436757E-09
C1 3 4 0.000012
Rpar 3 4 416666.666666667
.ends 870056174002_12uF
*******
.subckt 870056175003_22uF 1 2
Rser 1 3 0.0117190140844
Lser 2 4 5.170360925E-09
C1 3 4 0.000022
Rpar 3 4 227272.727272727
.ends 870056175003_22uF
*******
.subckt 870056175004_27uF 1 2
Rser 1 3 0.00869896893708
Lser 2 4 6.292043137E-09
C1 3 4 0.000027
Rpar 3 4 185185.185185185
.ends 870056175004_27uF
*******
.subckt 870056175005_33uF 1 2
Rser 1 3 0.010709292404
Lser 2 4 6.327349697E-09
C1 3 4 0.000033
Rpar 3 4 151515.151515152
.ends 870056175005_33uF
*******
