**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ASNP
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 865250140001_10uF 1 2
Rser 1 3 2.80207723226
Lser 2 4 8.79230402E-10
C1 3 4 0.00001
Rpar 3 4 2100000
.ends 865250140001_10uF
*******
.subckt 865250140002_22uF 1 2
Rser 1 3 2.79274851491
Lser 2 4 9.31010869E-10
C1 3 4 0.000022
Rpar 3 4 2100000
.ends 865250140002_22uF
*******
.subckt 865250142003_33uF 1 2
Rser 1 3 1.56920817768
Lser 2 4 2.849371314E-09
C1 3 4 0.000033
Rpar 3 4 2100000
.ends 865250142003_33uF
*******
.subckt 865250143004_47uF 1 2
Rser 1 3 1.17987154159
Lser 2 4 3.757449668E-09
C1 3 4 0.000047
Rpar 3 4 2100000
.ends 865250143004_47uF
*******
.subckt 865250145005_100uF 1 2
Rser 1 3 0.570596523699
Lser 2 4 4.427067613E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865250145005_100uF
*******
.subckt 865250149006_100uF 1 2
Rser 1 3 0.54
Lser 2 4 0.00000000325
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865250149006_100uF
*******
.subckt 865250153007_220uF 1 2
Rser 1 3 0.24
Lser 2 4 0.0000000031
C1 3 4 0.00022
Rpar 3 4 454545.454545454
.ends 865250153007_220uF
*******
.subckt 865250153008_330uF 1 2
Rser 1 3 0.245
Lser 2 4 0.0000000033
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865250153008_330uF
*******
.subckt 865250157009_470uF 1 2
Rser 1 3 0.155
Lser 2 4 0.0000000038
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 865250157009_470uF
*******
.subckt 865250157010_560uF 1 2
Rser 1 3 0.134
Lser 2 4 0.0000000042
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 865250157010_560uF
*******
.subckt 865250240001_10uF 1 2
Rser 1 3 1.93839512911
Lser 2 4 8.46868376E-10
C1 3 4 0.00001
Rpar 3 4 3333333.33333333
.ends 865250240001_10uF
*******
.subckt 865250242002_22uF 1 2
Rser 1 3 1.88026088686
Lser 2 4 2.596205262E-09
C1 3 4 0.000022
Rpar 3 4 3333333.33333333
.ends 865250242002_22uF
*******
.subckt 865250243003_33uF 1 2
Rser 1 3 1.24406533829
Lser 2 4 3.172719202E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865250243003_33uF
*******
.subckt 865250243004_47uF 1 2
Rser 1 3 1.24014138823
Lser 2 4 3.438243393E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865250243004_47uF
*******
.subckt 865250245005_100uF 1 2
Rser 1 3 0.405
Lser 2 4 0.000000000085
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865250245005_100uF
*******
.subckt 865250249006_100uF 1 2
Rser 1 3 0.545
Lser 2 4 0.00000000011
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865250249006_100uF
*******
.subckt 865250253007_220uF 1 2
Rser 1 3 0.24
Lser 2 4 0.0000000031
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865250253007_220uF
*******
.subckt 865250257008_330uF 1 2
Rser 1 3 0.155
Lser 2 4 0.0000000039
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 865250257008_330uF
*******
.subckt 865250340001_3.3uF 1 2
Rser 1 3 2.72046865757
Lser 2 4 7.96640782E-10
C1 3 4 0.0000033
Rpar 3 4 5333333.33333333
.ends 865250340001_3.3uF
*******
.subckt 865250340002_4.7uF 1 2
Rser 1 3 2.70410325988
Lser 2 4 1.388914622E-09
C1 3 4 0.0000047
Rpar 3 4 5333333.33333333
.ends 865250340002_4.7uF
*******
.subckt 865250340003_10uF 1 2
Rser 1 3 2.79476639021
Lser 2 4 1.643322931E-09
C1 3 4 0.00001
Rpar 3 4 5333333.33333333
.ends 865250340003_10uF
*******
.subckt 865250342004_22uF 1 2
Rser 1 3 1.5892159717
Lser 2 4 2.808957253E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865250342004_22uF
*******
.subckt 865250343005_33uF 1 2
Rser 1 3 1.58307606967
Lser 2 4 2.557750523E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865250343005_33uF
*******
.subckt 865250345006_47uF 1 2
Rser 1 3 0.784419193802
Lser 2 4 4.021731661E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865250345006_47uF
*******
.subckt 865250349007_47uF 1 2
Rser 1 3 0.763104389579
Lser 2 4 5.643364285E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865250349007_47uF
*******
.subckt 865250353008_100uF 1 2
Rser 1 3 0.346451201971
Lser 2 4 5.406836275E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865250353008_100uF
*******
.subckt 865250357009_220uF 1 2
Rser 1 3 0.148
Lser 2 4 0.0000000038
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 865250357009_220uF
*******
.subckt 865250440001_3.3uF 1 2
Rser 1 3 2.6398298091
Lser 2 4 9.96006788E-10
C1 3 4 0.0000033
Rpar 3 4 8333333.33333333
.ends 865250440001_3.3uF
*******
.subckt 865250440002_4.7uF 1 2
Rser 1 3 0.743400767868
Lser 2 4 4.268578394E-09
C1 3 4 0.0000047
Rpar 3 4 8333333.33333333
.ends 865250440002_4.7uF
*******
.subckt 865250442003_10uF 1 2
Rser 1 3 1.96914120053
Lser 2 4 2.355585585E-09
C1 3 4 0.00001
Rpar 3 4 8333333.33333333
.ends 865250442003_10uF
*******
.subckt 865250443004_22uF 1 2
Rser 1 3 1.14232876316
Lser 2 4 3.242713193E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865250443004_22uF
*******
.subckt 865250445005_33uF 1 2
Rser 1 3 0.804567270713
Lser 2 4 3.984118565E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865250445005_33uF
*******
.subckt 865250445007_47uF 1 2
Rser 1 3 0.791976036976
Lser 2 4 4.103503648E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865250445007_47uF
*******
.subckt 865250449006_33uF 1 2
Rser 1 3 0.858951290374
Lser 2 4 5.504779605E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865250449006_33uF
*******
.subckt 865250449008_47uF 1 2
Rser 1 3 1.09847379321
Lser 2 4 5.153002329E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865250449008_47uF
*******
.subckt 865250453009_100uF 1 2
Rser 1 3 0.365423369804
Lser 2 4 5.514284288E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 865250453009_100uF
*******
.subckt 865250540001_2.2uF 1 2
Rser 1 3 1.5
Lser 2 4 0.00000000000055
C1 3 4 0.0000022
Rpar 3 4 11666666.6666667
.ends 865250540001_2.2uF
*******
.subckt 865250540002_3.3uF 1 2
Rser 1 3 1.45
Lser 2 4 0.0000000000011
C1 3 4 0.0000033
Rpar 3 4 11666666.6666667
.ends 865250540002_3.3uF
*******
.subckt 865250540003_4.7uF 1 2
Rser 1 3 1.52
Lser 2 4 0.000000000001
C1 3 4 0.0000047
Rpar 3 4 11666666.6666667
.ends 865250540003_4.7uF
*******
.subckt 865250543004_10uF 1 2
Rser 1 3 1.15
Lser 2 4 0.000000000003
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865250543004_10uF
*******
.subckt 865250543005_22uF 1 2
Rser 1 3 1.29141365525
Lser 2 4 3.667878968E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545454
.ends 865250543005_22uF
*******
.subckt 865250553006_33uF 1 2
Rser 1 3 0.407511361224
Lser 2 4 5.304821546E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865250553006_33uF
*******
.subckt 865250553007_47uF 1 2
Rser 1 3 0.41010959413
Lser 2 4 5.052293425E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865250553007_47uF
*******
.subckt 865250640001_100nF 1 2
Rser 1 3 3.01499141338
Lser 2 4 1.697119497E-09
C1 3 4 0.0000001
Rpar 3 4 16666666.6666667
.ends 865250640001_100nF
*******
.subckt 865250640002_220nF 1 2
Rser 1 3 2.65882240175
Lser 2 4 1.420593501E-09
C1 3 4 0.00000022
Rpar 3 4 16666666.6666667
.ends 865250640002_220nF
*******
.subckt 865250640003_330nF 1 2
Rser 1 3 2.87397913513
Lser 2 4 1.742625339E-09
C1 3 4 0.00000033
Rpar 3 4 16666666.6666667
.ends 865250640003_330nF
*******
.subckt 865250640004_470nF 1 2
Rser 1 3 3.05159450863
Lser 2 4 1.740250613E-09
C1 3 4 0.00000047
Rpar 3 4 16666666.6666667
.ends 865250640004_470nF
*******
.subckt 865250640005_1uF 1 2
Rser 1 3 2.13099155466
Lser 2 4 5.6577995E-10
C1 3 4 0.000001
Rpar 3 4 16666666.6666667
.ends 865250640005_1uF
*******
.subckt 865250640006_2.2uF 1 2
Rser 1 3 2.5892374066
Lser 2 4 4.29438408E-10
C1 3 4 0.0000022
Rpar 3 4 16666666.6666667
.ends 865250640006_2.2uF
*******
.subckt 865250640007_3.3uF 1 2
Rser 1 3 2.36301447742
Lser 2 4 4.29438408E-10
C1 3 4 0.0000033
Rpar 3 4 16666666.6666667
.ends 865250640007_3.3uF
*******
.subckt 865250642008_4.7uF 1 2
Rser 1 3 2.4438319353
Lser 2 4 1.404618845E-09
C1 3 4 0.0000047
Rpar 3 4 16666666.6666667
.ends 865250642008_4.7uF
*******
.subckt 865250643009_10uF 1 2
Rser 1 3 1.86400650101
Lser 2 4 3.256825695E-09
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 865250643009_10uF
*******
.subckt 865250653010_22uF 1 2
Rser 1 3 0.477761621019
Lser 2 4 4.997014336E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 865250653010_22uF
*******
.subckt 865250657011_33uF 1 2
Rser 1 3 0.165
Lser 2 4 0.0000000009
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 865250657011_33uF
*******
.subckt 865250657012_47uF 1 2
Rser 1 3 0.165
Lser 2 4 0.0000000009
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 865250657012_47uF
*******
