**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Rod Core Inductor SMT
* Matchcode:             WE-RCIS
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/8/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 7847227010_1u 1 2
Rp 1 2 4761
Cp 1 2 0.96078p
Rs 1 N3 0.002
L1 N3 2 0.615082u
.ends 7847227010_1u
*******
.subckt 7847227027_2.72u 1 2
Rp 1 2 11385
Cp 1 2 1.139p
Rs 1 N3 0.0064
L1 N3 2 1.547u
.ends 7847227027_2.72u
*******
.subckt 7847229020_1.96u 1 2
Rp 1 2 10064
Cp 1 2 1.214p
Rs 1 N3 0.0024
L1 N3 2 1.147u
.ends 7847229020_1.96u
*******
.subckt 7847232045_4.45u 1 2
Rp 1 2 3427
Cp 1 2 4.56p
Rs 1 N3 0.0038
L1 N3 2 3.237u
.ends 7847232045_4.45u
*******
