**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Multilayer Ceramic Chip Capacitors
* Matchcode:             WCAP-CSRF
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0201_885392004001_0.2pF 1 2
Rser 1 3 0.601
Lser 2 4 0.000000000325
C1 3 4 0.00000000000025
Rpar 3 4 10000000000
.ends 0201_885392004001_0.2pF
*******
.subckt 0201_885392004002_1pF 1 2
Rser 1 3 0.409
Lser 2 4 0.000000000365
C1 3 4 0.00000000000105
Rpar 3 4 10000000000
.ends 0201_885392004002_1pF
*******
.subckt 0201_885392004003_1.2pF 1 2
Rser 1 3 0.386
Lser 2 4 0.000000000395
C1 3 4 0.00000000000126
Rpar 3 4 10000000000
.ends 0201_885392004003_1.2pF
*******
.subckt 0201_885392004004_1.5pF 1 2
Rser 1 3 0.368
Lser 2 4 0.00000000039
C1 3 4 0.00000000000157
Rpar 3 4 10000000000
.ends 0201_885392004004_1.5pF
*******
.subckt 0201_885392004005_2.2pF 1 2
Rser 1 3 0.335
Lser 2 4 0.00000000037
C1 3 4 0.00000000000227
Rpar 3 4 10000000000
.ends 0201_885392004005_2.2pF
*******
.subckt 0201_885392004006_2.7pF 1 2
Rser 1 3 0.285
Lser 2 4 0.000000000345
C1 3 4 0.00000000000276
Rpar 3 4 10000000000
.ends 0201_885392004006_2.7pF
*******
.subckt 0201_885392004007_3.3pF 1 2
Rser 1 3 0.256
Lser 2 4 0.00000000039
C1 3 4 0.00000000000338
Rpar 3 4 10000000000
.ends 0201_885392004007_3.3pF
*******
.subckt 0201_885392004008_4.7pF 1 2
Rser 1 3 0.203
Lser 2 4 0.00000000038
C1 3 4 0.00000000000478
Rpar 3 4 10000000000
.ends 0201_885392004008_4.7pF
*******
.subckt 0201_885392004009_5.6pF 1 2
Rser 1 3 0.193
Lser 2 4 0.00000000039
C1 3 4 0.00000000000574
Rpar 3 4 10000000000
.ends 0201_885392004009_5.6pF
*******
.subckt 0201_885392004010_9pF 1 2
Rser 1 3 0.155
Lser 2 4 0.0000000004
C1 3 4 0.00000000000916
Rpar 3 4 10000000000
.ends 0201_885392004010_9pF
*******
.subckt 0201_885392004011_33pF 1 2
Rser 1 3 0.0858
Lser 2 4 0.00000000037
C1 3 4 0.0000000000333
Rpar 3 4 10000000000
.ends 0201_885392004011_33pF
*******
.subckt 0402_885392005001_0.3pF 1 2
Rser 1 3 0.736
Lser 2 4 0.0000000003
C1 3 4 0.000000000000365
Rpar 3 4 10000000000
.ends 0402_885392005001_0.3pF
*******
.subckt 0402_885392005002_0.4pF 1 2
Rser 1 3 0.693
Lser 2 4 0.00000000034
C1 3 4 0.000000000000467
Rpar 3 4 10000000000
.ends 0402_885392005002_0.4pF
*******
.subckt 0402_885392005003_0.4pF 1 2
Rser 1 3 0.693
Lser 2 4 0.00000000034
C1 3 4 0.000000000000467
Rpar 3 4 10000000000
.ends 0402_885392005003_0.4pF
*******
.subckt 0402_885392005004_0.5pF 1 2
Rser 1 3 0.634
Lser 2 4 0.00000000035
C1 3 4 0.000000000000571
Rpar 3 4 10000000000
.ends 0402_885392005004_0.5pF
*******
.subckt 0402_885392005005_1pF 1 2
Rser 1 3 0.506
Lser 2 4 0.0000000005
C1 3 4 0.00000000000108
Rpar 3 4 10000000000
.ends 0402_885392005005_1pF
*******
.subckt 0402_885392005006_1pF 1 2
Rser 1 3 0.506
Lser 2 4 0.0000000005
C1 3 4 0.00000000000108
Rpar 3 4 10000000000
.ends 0402_885392005006_1pF
*******
.subckt 0402_885392005007_1.5pF 1 2
Rser 1 3 0.473
Lser 2 4 0.00000000045
C1 3 4 0.00000000000161
Rpar 3 4 10000000000
.ends 0402_885392005007_1.5pF
*******
.subckt 0402_885392005008_1.8pF 1 2
Rser 1 3 0.443
Lser 2 4 0.00000000047
C1 3 4 0.00000000000188
Rpar 3 4 10000000000
.ends 0402_885392005008_1.8pF
*******
.subckt 0402_885392005009_2.3pF 1 2
Rser 1 3 0.363
Lser 2 4 0.0000000004
C1 3 4 0.00000000000242
Rpar 3 4 10000000000
.ends 0402_885392005009_2.3pF
*******
.subckt 0402_885392005010_3pF 1 2
Rser 1 3 0.273
Lser 2 4 0.0000000004
C1 3 4 0.00000000000308
Rpar 3 4 10000000000
.ends 0402_885392005010_3pF
*******
.subckt 0402_885392005011_3.3pF 1 2
Rser 1 3 0.52
Lser 2 4 0.0000000004
C1 3 4 0.00000000000339
Rpar 3 4 10000000000
.ends 0402_885392005011_3.3pF
*******
.subckt 0402_885392005012_4.7pF 1 2
Rser 1 3 0.21
Lser 2 4 0.00000000044
C1 3 4 0.00000000000481
Rpar 3 4 10000000000
.ends 0402_885392005012_4.7pF
*******
.subckt 0402_885392005013_5.6pF 1 2
Rser 1 3 0.92
Lser 2 4 0.00000000044
C1 3 4 0.00000000000566
Rpar 3 4 10000000000
.ends 0402_885392005013_5.6pF
*******
.subckt 0402_885392005014_9pF 1 2
Rser 1 3 0.164
Lser 2 4 0.000000000507
C1 3 4 0.00000000000906
Rpar 3 4 10000000000
.ends 0402_885392005014_9pF
*******
