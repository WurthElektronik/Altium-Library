**************************************************
* Manufacturer:           Würth Elektronik
* Kinds:                  SMT Mono-color Chip LED Diffused
* Matchcode:              WL-SMCD
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2024-01-26
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2024 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0603_150060AS55040 1 2
D1 1 2 SMCD
.MODEL SMCD D
+ IS=179.05E-12
+ N=4.1622
+ RS=.56312
+ IKF=81.248
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
*****************************
.subckt 0603_150060BS55040 1 2
D1 1 2 SMCD
.MODEL SMCD D
+ IS=11.416E-15
+ N=3.7886
+ RS=1.4842
+ IKF=213.88E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
*****************************
.subckt 0603_150060GS55040 1 2
D1 1 2 SMCD
.MODEL SMCD D
+ IS=406.49E-12
+ N=4.8627
+ RS=4.1370
+ IKF=13.914E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
*****************************
.subckt 0603_150060RS55040 1 2
D1 1 2 SMCD
.MODEL SMCD D
+ IS=153.31E-12
+ N=4.1406
+ RS=1.0267
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
*****************************
.subckt 0603_150060SS55040 1 2
D1 1 2 SMCD
.MODEL SMCD D
+ IS=153.31E-12
+ N=4.1406
+ RS=1.0267
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
*****************************
.subckt 0603_150060YS55040 1 2
D1 1 2 SMCD
.MODEL SMCD D
+ IS=135.21E-15
+ N=2.0992
+ RS=1.0413
+ IKF=173.47E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
*****************************
.subckt 0603_150060VS55040 1 2
D1 1 2 SMCD
.MODEL SMCD D
+ IS=135.21E-15
+ N=2.0992
+ RS=1.0413
+ IKF=173.47E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
+ TT=5.0000E-9
.ends
*****************************

