**************************************************
* Manufacturer:          W�rth Elektronik
* Kinds:                 SMT Power Inductor
* Matchcode:             WE-MAIA
* Library Type:          LTspice
* Version:               rev24a
* Created/modified by:   Ella
* Date and Time:         2024/09/13
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2024 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 2512_784383240047_0.47u 1 2
Rp 1 2 1038.4604951
Cp 1 2 2.9596p
Rs 1 N3 0.03
L1 N3 2 0.39u
.ends 2512_784383240047_0.47u
*******
.subckt 2512_784383240056_0.56u 1 2
Rp 1 2 1377.704037902
Cp 1 2 3.265353363p
Rs 1 N3 0.037
L1 N3 2 0.53u
.ends 2512_784383240056_0.56u
*******
.subckt 2512_784383240068_0.68u 1 2
Rp 1 2 1711.275912736
Cp 1 2 3.4284831524p
Rs 1 N3 0.045
L1 N3 2 0.66u
.ends 2512_784383240068_0.68u
*******
.subckt 2512_78438324010_1u 1 2
Rp 1 2 2168.089901022
Cp 1 2 3.75836481733333p
Rs 1 N3 0.049
L1 N3 2 0.93u
.ends 2512_78438324010_1u
*******
.subckt 2512_78438324012_1.2u 1 2
Rp 1 2 2597.705977778
Cp 1 2 3.9005958574p
Rs 1 N3 0.067
L1 N3 2 1.07u
.ends 2512_78438324012_1.2u
*******
.subckt 2512_78438324015_1.5u 1 2
Rp 1 2 3445.783694548
Cp 1 2 4.425720698p
Rs 1 N3 0.082
L1 N3 2 1.54u
.ends 2512_78438324015_1.5u
*******
.subckt 2512_78438324022_2.2u 1 2
Rp 1 2 4211.982563034
Cp 1 2 4.0585787336p
Rs 1 N3 0.123
L1 N3 2 1.87u
.ends 2512_78438324022_2.2u
*******
.subckt 2512_78438324033_3.3u 1 2
Rp 1 2 7042.196136376
Cp 1 2 4.3926298308p
Rs 1 N3 0.226
L1 N3 2 3.25u
.ends 2512_78438324033_3.3u
*******
.subckt 2512_78438324047_4.7u 1 2
Rp 1 2 9138.238352662
Cp 1 2 4.3223636442p
Rs 1 N3 0.3
L1 N3 2 4.48u
.ends 2512_78438324047_4.7u
*******
.subckt 2512_78438324056_5.6u 1 2
Rp 1 2 10933.60876782
Cp 1 2 5.1948829364p
Rs 1 N3 0.405
L1 N3 2 5.69u
.ends 2512_78438324056_5.6u
*******
.subckt 2512_78438324068_6.8u 1 2
Rp 1 2 12309.69262034
Cp 1 2 4.9992358046p
Rs 1 N3 0.56
L1 N3 2 6.69u
.ends 2512_78438324068_6.8u
*******
.subckt 2512_78438324082_8.2u 1 2
Rp 1 2 14021.69415194
Cp 1 2 5.0174407148p
Rs 1 N3 0.63
L1 N3 2 7.88u
.ends 2512_78438324082_8.2u
*******
.subckt 2506_784383210047_0.47u 1 2
Rp 1 2 1358.795
Cp 1 2 2.20133333333333p
Rs 1 N3 0.076
L1 N3 2 0.49u
.ends 2506_784383210047_0.47u
*******
.subckt 2506_78438321010_1u 1 2
Rp 1 2 2580.266667
Cp 1 2 2.89383333333333p
Rs 1 N3 0.163
L1 N3 2 1.09u
.ends 2506_78438321010_1u
*******
.subckt 2508_784383220047_0.47u 1 2
Rp 1 2 1328.67
Cp 1 2 2.363p
Rs 1 N3 0.07
L1 N3 2 0.48u
.ends 2508_784383220047_0.47u
*******
.subckt 2508_78438322010_1u 1 2
Rp 1 2 2287
Cp 1 2 2.785p
Rs 1 N3 0.107
L1 N3 2 0.93u
.ends 2508_78438322010_1u
*******
.subckt 2508_78438322022_2.2u 1 2
Rp 1 2 5454.6
Cp 1 2 3.2106p
Rs 1 N3 0.252
L1 N3 2 2.4u
.ends 2508_78438322022_2.2u
*******
.subckt 2510_784383230033_0.33u 1 2
Rp 1 2 759.73
Cp 1 2 2.78833333333333p
Rs 1 N3 0.029
L1 N3 2 0.28u
.ends 2510_784383230033_0.33u
*******
.subckt 2510_784383230047_0.47u 1 2
Rp 1 2 807.55
Cp 1 2 2.235p
Rs 1 N3 0.037
L1 N3 2 0.44u
.ends 2510_784383230047_0.47u
*******
.subckt 2510_784383230068_0.68u 1 2
Rp 1 2 1052.9
Cp 1 2 2.57566666666667p
Rs 1 N3 0.046
L1 N3 2 0.62u
.ends 2510_784383230068_0.68u
*******
.subckt 2510_784383230082_0.82u 1 2
Rp 1 2 1712.77
Cp 1 2 3.18373333333333p
Rs 1 N3 0.053
L1 N3 2 0.77u
.ends 2510_784383230082_0.82u
*******
.subckt 2510_78438323010_1u 1 2
Rp 1 2 2155.33
Cp 1 2 3.992p
Rs 1 N3 0.063
L1 N3 2 1.01u
.ends 2510_78438323010_1u
*******
.subckt 2510_78438323012_1.2u 1 2
Rp 1 2 2888.67
Cp 1 2 3.38366666666667p
Rs 1 N3 0.082
L1 N3 2 1.2u
.ends 2510_78438323012_1.2u
*******
.subckt 2510_78438323015_1.5u 1 2
Rp 1 2 3356.67
Cp 1 2 3.701p
Rs 1 N3 0.092
L1 N3 2 1.41u
.ends 2510_78438323015_1.5u
*******
.subckt 2510_78438323022_2.2u 1 2
Rp 1 2 2863
Cp 1 2 2.63366666666667p
Rs 1 N3 0.147
L1 N3 2 2.3u
.ends 2510_78438323022_2.2u
*******
.subckt 2510_78438323033_3.3u 1 2
Rp 1 2 5818.67
Cp 1 2 3.66p
Rs 1 N3 0.22
L1 N3 2 3.01u
.ends 2510_78438323033_3.3u
*******
.subckt 2510_78438323047_4.7u 1 2
Rp 1 2 8723.67
Cp 1 2 4.55633333333333p
Rs 1 N3 0.338
L1 N3 2 4.61u
.ends 2510_78438323047_4.7u
*******
.subckt 2510_78438323068_6.8u 1 2
Rp 1 2 12938.33
Cp 1 2 3.90866666666667p
Rs 1 N3 0.563
L1 N3 2 6.51u
.ends 2510_78438323068_6.8u
*******
.subckt 2510_78438323082_8.2u 1 2
Rp 1 2 14641.63
Cp 1 2 4.42933333333333p
Rs 1 N3 0.646
L1 N3 2 8.12u
.ends 2510_78438323082_8.2u
*******
.subckt 2510_78438323100_10u 1 2
Rp 1 2 17001.67
Cp 1 2 4.38766666666667p
Rs 1 N3 0.733
L1 N3 2 9.66u
.ends 2510_78438323100_10u
*******
.subckt 2512_78438324100_10u 1 2
Rp 1 2 13964.0031297
Cp 1 2 4.94140041425p
Rs 1 N3 0.68
L1 N3 2 8.13u
.ends 2512_78438324100_10u
*******
.subckt 3010_78438333022_2.2u 1 2
Rp 1 2 5803.666667
Cp 1 2 4.724p
Rs 1 N3 0.15
L1 N3 2 2.1u
.ends 3010_78438333022_2.2u
*******
.subckt 3010_78438333033_3.3u 1 2
Rp 1 2 8309.333333
Cp 1 2 5.34966666666667p
Rs 1 N3 0.232
L1 N3 2 3.09u
.ends 3010_78438333033_3.3u
*******
.subckt 3010_78438333047_4.7u 1 2
Rp 1 2 8564.333333
Cp 1 2 5.27933333333333p
Rs 1 N3 0.356
L1 N3 2 4.45u
.ends 3010_78438333047_4.7u
*******
.subckt 3012_784383340033_0.33u 1 2
Rp 1 2 821.2233333
Cp 1 2 4.27333333333333p
Rs 1 N3 0.019
L1 N3 2 0.29u
.ends 3012_784383340033_0.33u
*******
.subckt 3012_784383340047_0.47u 1 2
Rp 1 2 1173.333333
Cp 1 2 4.55666666666667p
Rs 1 N3 0.022
L1 N3 2 0.4u
.ends 3012_784383340047_0.47u
*******
.subckt 3012_784383340056_0.56u 1 2
Rp 1 2 1565
Cp 1 2 3.79066666666667p
Rs 1 N3 0.029
L1 N3 2 0.57u
.ends 3012_784383340056_0.56u
*******
.subckt 3012_784383340068_0.68u 1 2
Rp 1 2 1736.666667
Cp 1 2 3.80966666666667p
Rs 1 N3 0.036
L1 N3 2 0.65u
.ends 3012_784383340068_0.68u
*******
.subckt 3012_78438334010_1u 1 2
Rp 1 2 2542.333333
Cp 1 2 4.17533333333333p
Rs 1 N3 0.0421
L1 N3 2 1.08u
.ends 3012_78438334010_1u
*******
.subckt 3012_78438334012_1.2u 1 2
Rp 1 2 3020.5
Cp 1 2 4.95453333333333p
Rs 1 N3 0.055
L1 N3 2 1.22u
.ends 3012_78438334012_1.2u
*******
.subckt 3012_78438334015_1.5u 1 2
Rp 1 2 3865
Cp 1 2 4.74866666666667p
Rs 1 N3 0.08
L1 N3 2 1.5u
.ends 3012_78438334015_1.5u
*******
.subckt 3012_78438334022_2.2u 1 2
Rp 1 2 4887.666667
Cp 1 2 5.10166666666667p
Rs 1 N3 0.1
L1 N3 2 2.04u
.ends 3012_78438334022_2.2u
*******
.subckt 3012_78438334033_3.3u 1 2
Rp 1 2 7481
Cp 1 2 6.07033333333333p
Rs 1 N3 0.1563
L1 N3 2 3.26u
.ends 3012_78438334033_3.3u
*******
.subckt 3012_78438334047_4.7u 1 2
Rp 1 2 9053.666667
Cp 1 2 5.97833333333333p
Rs 1 N3 0.2677
L1 N3 2 4.38u
.ends 3012_78438334047_4.7u
*******
.subckt 3012_78438334056_5.6u 1 2
Rp 1 2 10141
Cp 1 2 5.743p
Rs 1 N3 0.3383
L1 N3 2 5.5u
.ends 3012_78438334056_5.6u
*******
.subckt 3012_78438334068_6.8u 1 2
Rp 1 2 11556.33333
Cp 1 2 6.09933333333333p
Rs 1 N3 0.3682
L1 N3 2 5.99u
.ends 3012_78438334068_6.8u
*******
.subckt 3015_784383350047_0.47u 1 2
Rp 1 2 1058.19523333333
Cp 1 2 4.85417386666667p
Rs 1 N3 0.02
L1 N3 2 0.45u
.ends 3015_784383350047_0.47u
*******
.subckt 3015_784383350068_0.68u 1 2
Rp 1 2 1639.15646368427
Cp 1 2 4.395p
Rs 1 N3 0.025
L1 N3 2 0.51u
.ends 3015_784383350068_0.68u
*******
.subckt 3015_784383350082_0.82u 1 2
Rp 1 2 2232.88336666667
Cp 1 2 4.5684805p
Rs 1 N3 0.03
L1 N3 2 0.75u
.ends 3015_784383350082_0.82u
*******
.subckt 3015_78438335010_1u 1 2
Rp 1 2 2039.333333
Cp 1 2 4.95603333333333p
Rs 1 N3 0.039
L1 N3 2 1.02u
.ends 3015_78438335010_1u
*******
.subckt 3015_78438335022_2.2u 1 2
Rp 1 2 4443
Cp 1 2 5.69266666666667p
Rs 1 N3 0.094
L1 N3 2 1.98u
.ends 3015_78438335022_2.2u
*******
.subckt 3015_78438335033_3.3u 1 2
Rp 1 2 6061
Cp 1 2 6.48433333333333p
Rs 1 N3 0.114
L1 N3 2 3.13u
.ends 3015_78438335033_3.3u
*******
.subckt 3015_78438335047_4.7u 1 2
Rp 1 2 8005.666667
Cp 1 2 6.65533333333333p
Rs 1 N3 0.141
L1 N3 2 4.26u
.ends 3015_78438335047_4.7u
*******
.subckt 3015_78438335068_6.8u 1 2
Rp 1 2 10791.66667
Cp 1 2 7.02333333333333p
Rs 1 N3 0.25
L1 N3 2 6.25u
.ends 3015_78438335068_6.8u
*******
.subckt 3015_78438335100_10u 1 2
Rp 1 2 15109.66667
Cp 1 2 6.18366666666667p
Rs 1 N3 0.446
L1 N3 2 9.46u
.ends 3015_78438335100_10u
*******
.subckt 3015_78438335150_15u 1 2
Rp 1 2 21284.66667
Cp 1 2 5.87033333333333p
Rs 1 N3 0.72
L1 N3 2 14.1u
.ends 3015_78438335150_15u
*******
.subckt 3015_78438335220_22u 1 2
Rp 1 2 29029
Cp 1 2 6.34333333333333p
Rs 1 N3 0.94
L1 N3 2 19.78u
.ends 3015_78438335220_22u
*******
.subckt 3015_78438335330_33u 1 2
Rp 1 2 33248.33333
Cp 1 2 6.99333333333333p
Rs 1 N3 1.21
L1 N3 2 29.66u
.ends 3015_78438335330_33u
*******
.subckt 3015_78438335470_47u 1 2
Rp 1 2 42066.66667
Cp 1 2 7.59833333333333p
Rs 1 N3 2.09
L1 N3 2 46.1u
.ends 3015_78438335470_47u
*******
.subckt 3020_784383360033_0.33u 1 2
Rp 1 2 725.017800117
Cp 1 2 4.2139562698p
Rs 1 N3 0.014
L1 N3 2 0.31u
.ends 3020_784383360033_0.33u
*******
.subckt 3020_784383360047_0.47u 1 2
Rp 1 2 1054.617100708
Cp 1 2 5.3828993388p
Rs 1 N3 0.018
L1 N3 2 0.46u
.ends 3020_784383360047_0.47u
*******
.subckt 3020_784383360068_0.68u 1 2
Rp 1 2 1402.486795318
Cp 1 2 5.6011470144p
Rs 1 N3 0.022
L1 N3 2 0.65u
.ends 3020_784383360068_0.68u
*******
.subckt 3020_78438336010_1u 1 2
Rp 1 2 1905.123596372
Cp 1 2 5.8797906294p
Rs 1 N3 0.026
L1 N3 2 0.95u
.ends 3020_78438336010_1u
*******
.subckt 3020_78438336012_1.2u 1 2
Rp 1 2 2327.00997736
Cp 1 2 6.4008161236p
Rs 1 N3 0.03
L1 N3 2 1.18u
.ends 3020_78438336012_1.2u
*******
.subckt 3020_78438336015_1.5u 1 2
Rp 1 2 2879.288208634
Cp 1 2 6.5500806518p
Rs 1 N3 0.033
L1 N3 2 1.46u
.ends 3020_78438336015_1.5u
*******
.subckt 3020_78438336022_2.2u 1 2
Rp 1 2 4907.58956685
Cp 1 2 6.44236118p
Rs 1 N3 0.067
L1 N3 2 2.22u
.ends 3020_78438336022_2.2u
*******
.subckt 3020_78438336033_3.3u 1 2
Rp 1 2 6097.32637741
Cp 1 2 5.7471916388p
Rs 1 N3 0.099
L1 N3 2 2.92u
.ends 3020_78438336033_3.3u
*******
.subckt 3020_78438336047_4.7u 1 2
Rp 1 2 8959.521080854
Cp 1 2 6.4455729074p
Rs 1 N3 0.137
L1 N3 2 4.52u
.ends 3020_78438336047_4.7u
*******
.subckt 3020_78438336068_6.8u 1 2
Rp 1 2 9175.279119816
Cp 1 2 8.1999260564p
Rs 1 N3 0.168
L1 N3 2 6.23u
.ends 3020_78438336068_6.8u
*******
.subckt 3020_78438336100_10u 1 2
Rp 1 2 14215.45725152
Cp 1 2 8.016436544p
Rs 1 N3 0.28
L1 N3 2 9.07u
.ends 3020_78438336100_10u
*******
.subckt 4020_784383560033_0.33u 1 2
Rp 1 2 710
Cp 1 2 5.49p
Rs 1 N3 0.006
L1 N3 2 0.32u
.ends 4020_784383560033_0.33u
*******
.subckt 4020_784383560056_0.56u 1 2
Rp 1 2 1091
Cp 1 2 5.821p
Rs 1 N3 0.007
L1 N3 2 0.49u
.ends 4020_784383560056_0.56u
*******
.subckt 4020_784383560068_0.68u 1 2
Rp 1 2 1329
Cp 1 2 7.075p
Rs 1 N3 0.0075
L1 N3 2 0.63u
.ends 4020_784383560068_0.68u
*******
.subckt 4020_78438356010_1u 1 2
Rp 1 2 2207
Cp 1 2 8.5p
Rs 1 N3 0.012
L1 N3 2 1.01u
.ends 4020_78438356010_1u
*******
.subckt 4020_78438356012_1.2u 1 2
Rp 1 2 2437
Cp 1 2 7.5p
Rs 1 N3 0.015
L1 N3 2 1.15u
.ends 4020_78438356012_1.2u
*******
.subckt 4020_78438356015_1.5u 1 2
Rp 1 2 2807
Cp 1 2 8.18p
Rs 1 N3 0.016
L1 N3 2 1.38u
.ends 4020_78438356015_1.5u
*******
.subckt 4020_78438356018_1.8u 1 2
Rp 1 2 3494
Cp 1 2 8.87p
Rs 1 N3 0.0245
L1 N3 2 1.79u
.ends 4020_78438356018_1.8u
*******
.subckt 4020_78438356022_2.2u 1 2
Rp 1 2 3998
Cp 1 2 9.56p
Rs 1 N3 0.029
L1 N3 2 2.18u
.ends 4020_78438356022_2.2u
*******
.subckt 4020_78438356033_3.3u 1 2
Rp 1 2 5464
Cp 1 2 12.635p
Rs 1 N3 0.0399
L1 N3 2 3.18u
.ends 4020_78438356033_3.3u
*******
.subckt 4020_78438356047_4.7u 1 2
Rp 1 2 7282
Cp 1 2 11.809p
Rs 1 N3 0.063
L1 N3 2 4.67u
.ends 4020_78438356047_4.7u
*******
.subckt 4020_78438356056_5.6u 1 2
Rp 1 2 8507
Cp 1 2 11.152p
Rs 1 N3 0.068
L1 N3 2 5.17u
.ends 4020_78438356056_5.6u
*******
.subckt 4030_78438357010_1u 1 2
Rp 1 2 2195
Cp 1 2 7.039p
Rs 1 N3 0.0116
L1 N3 2 0.95u
.ends 4030_78438357010_1u
*******
.subckt 4030_78438357012_1.2u 1 2
Rp 1 2 2666
Cp 1 2 7.978933146p
Rs 1 N3 0.0134
L1 N3 2 1.22u
.ends 4030_78438357012_1.2u
*******
.subckt 4030_78438357015_1.5u 1 2
Rp 1 2 3039
Cp 1 2 7.847855157p
Rs 1 N3 0.0171
L1 N3 2 1.37u
.ends 4030_78438357015_1.5u
*******
.subckt 4030_78438357018_1.8u 1 2
Rp 1 2 3649
Cp 1 2 8.081p
Rs 1 N3 0.018
L1 N3 2 1.7u
.ends 4030_78438357018_1.8u
*******
.subckt 4030_78438357022_2.2u 1 2
Rp 1 2 4556
Cp 1 2 9.489572495p
Rs 1 N3 0.022
L1 N3 2 2.11u
.ends 4030_78438357022_2.2u
*******
.subckt 4030_78438357033_3.3u 1 2
Rp 1 2 4719
Cp 1 2 11.849p
Rs 1 N3 0.029
L1 N3 2 3.236u
.ends 4030_78438357033_3.3u
*******
.subckt 4030_78438357047_4.7u 1 2
Rp 1 2 8253
Cp 1 2 10.011598369p
Rs 1 N3 0.0399
L1 N3 2 4.22u
.ends 4030_78438357047_4.7u
*******
.subckt 4030_78438357056_5.6u 1 2
Rp 1 2 9277
Cp 1 2 11.153505232p
Rs 1 N3 0.0465
L1 N3 2 5.7u
.ends 4030_78438357056_5.6u
*******
.subckt 4030_78438357068_6.8u 1 2
Rp 1 2 11078
Cp 1 2 10p
Rs 1 N3 0.0694
L1 N3 2 6.45u
.ends 4030_78438357068_6.8u
*******
.subckt 4030_78438357082_8.2u 1 2
Rp 1 2 12230
Cp 1 2 11.388p
Rs 1 N3 0.081
L1 N3 2 7.76u
.ends 4030_78438357082_8.2u
*******
.subckt 4030_78438357100_10u 1 2
Rp 1 2 13721
Cp 1 2 11.841p
Rs 1 N3 0.1008
L1 N3 2 9.47u
.ends 4030_78438357100_10u
*******
.subckt 1610_784383130033_0.33u 1 2
Rp 1 2 1175.839
Cp 1 2 1.6355p
Rs 1 N3 0.065
L1 N3 2 0.346u
.ends 1610_784383130033_0.33u
*******
.subckt 1610_784383130047_0.47u 1 2
Rp 1 2 1548.746
Cp 1 2 1.657p
Rs 1 N3 0.077
L1 N3 2 0.52u
.ends 1610_784383130047_0.47u
*******
.subckt 1610_784383130056_0.56u 1 2
Rp 1 2 1864.888
Cp 1 2 1.8707p
Rs 1 N3 0.09
L1 N3 2 0.58u
.ends 1610_784383130056_0.56u
*******
.subckt 1610_784383130068_0.68u 1 2
Rp 1 2 2230.246
Cp 1 2 1.9747p
Rs 1 N3 0.101
L1 N3 2 0.74u
.ends 1610_784383130068_0.68u
*******
.subckt 1610_784383130082_0.82u 1 2
Rp 1 2 2577.813
Cp 1 2 2.153p
Rs 1 N3 0.115
L1 N3 2 0.9u
.ends 1610_784383130082_0.82u
*******
.subckt 1610_78438313010_1u 1 2
Rp 1 2 3023.53
Cp 1 2 2.1174p
Rs 1 N3 0.127
L1 N3 2 0.99u
.ends 1610_78438313010_1u
*******
.subckt 1610_78438313012_1.2u 1 2
Rp 1 2 3481.561
Cp 1 2 2.0866p
Rs 1 N3 0.14
L1 N3 2 1.18u
.ends 1610_78438313012_1.2u
*******
.subckt 1610_78438313015_1.5u 1 2
Rp 1 2 4017.414
Cp 1 2 2.5328p
Rs 1 N3 0.189
L1 N3 2 1.46u
.ends 1610_78438313015_1.5u
*******
.subckt 1610_78438313022_2.2u 1 2
Rp 1 2 5651.21
Cp 1 2 2.5307p
Rs 1 N3 0.337
L1 N3 2 2.27u
.ends 1610_78438313022_2.2u
*******
.subckt 4020HT_784383560033HT_0.33u 1 2
Rp 1 2 713.426
Cp 1 2 7.731p
Rs 1 N3 0.0065
L1 N3 2 0.376u
.ends 4020HT_784383560033HT_0.33u
*******
.subckt 4020HT_784383560047HT_0.47u 1 2
Rp 1 2 970.242
Cp 1 2 8.284p
Rs 1 N3 0.007
L1 N3 2 0.485199u
.ends 4020HT_784383560047HT_0.47u
*******
.subckt 4020HT_784383560056HT_0.56u 1 2
Rp 1 2 1279
Cp 1 2 8.414p
Rs 1 N3 0.0075
L1 N3 2 0.603265u
.ends 4020HT_784383560056HT_0.56u
*******
.subckt 4020HT_784383560068HT_0.68u 1 2
Rp 1 2 1382
Cp 1 2 9.284p
Rs 1 N3 0.008
L1 N3 2 0.637919u
.ends 4020HT_784383560068HT_0.68u
*******
.subckt 4020HT_78438356010HT_1u 1 2
Rp 1 2 2276
Cp 1 2 10.825p
Rs 1 N3 0.0135
L1 N3 2 1.168u
.ends 4020HT_78438356010HT_1u
*******
.subckt 4020HT_78438356012HT_1.2u 1 2
Rp 1 2 2454
Cp 1 2 10.374p
Rs 1 N3 0.016
L1 N3 2 1.325u
.ends 4020HT_78438356012HT_1.2u
*******
.subckt 4020HT_78438356015HT_1.5u 1 2
Rp 1 2 2780
Cp 1 2 10.604p
Rs 1 N3 0.018
L1 N3 2 1.55u
.ends 4020HT_78438356015HT_1.5u
*******
.subckt 4020HT_78438356018HT_1.8u 1 2
Rp 1 2 3724
Cp 1 2 9.572p
Rs 1 N3 0.026
L1 N3 2 1.961u
.ends 4020HT_78438356018HT_1.8u
*******
.subckt 4020HT_78438356022HT_2.2u 1 2
Rp 1 2 4107
Cp 1 2 12.2p
Rs 1 N3 0.028
L1 N3 2 2.328u
.ends 4020HT_78438356022HT_2.2u
*******
.subckt 4020HT_78438356033HT_3.3u 1 2
Rp 1 2 6048
Cp 1 2 12.082p
Rs 1 N3 0.045
L1 N3 2 3.55u
.ends 4020HT_78438356033HT_3.3u
*******
.subckt 4020HT_78438356047HT_4.7u 1 2
Rp 1 2 7131
Cp 1 2 14.902p
Rs 1 N3 0.065
L1 N3 2 5.262u
.ends 4020HT_78438356047HT_4.7u
*******
.subckt 4020HT_78438356056HT_5.6u 1 2
Rp 1 2 7849
Cp 1 2 15.226p
Rs 1 N3 0.07
L1 N3 2 5.699u
.ends 4020HT_78438356056HT_5.6u
*******
.subckt 5020_784383660082_0.82u 1 2
Rp 1 2 1355
Cp 1 2 11.133p
Rs 1 N3 0.0083
L1 N3 2 0.796u
.ends 5020_784383660082_0.82u
*******
.subckt 5020_78438366010_1u 1 2
Rp 1 2 1863
Cp 1 2 11.252p
Rs 1 N3 0.0114
L1 N3 2 1.016u
.ends 5020_78438366010_1u
*******
.subckt 5020_78438366015_1.5u 1 2
Rp 1 2 2481
Cp 1 2 11.154p
Rs 1 N3 0.0185
L1 N3 2 1.618u
.ends 5020_78438366015_1.5u
*******
.subckt 5020_78438366022_2.2u 1 2
Rp 1 2 3190
Cp 1 2 12.557p
Rs 1 N3 0.0237
L1 N3 2 2.037u
.ends 5020_78438366022_2.2u
*******
.subckt 5020_78438366033_3.3u 1 2
Rp 1 2 4100
Cp 1 2 14.524p
Rs 1 N3 0.0334
L1 N3 2 3.202u
.ends 5020_78438366033_3.3u
*******
.subckt 5020_78438366047_4.7u 1 2
Rp 1 2 4923
Cp 1 2 14.429p
Rs 1 N3 0.0548
L1 N3 2 4.483u
.ends 5020_78438366047_4.7u
*******
.subckt 5030_78438367010_1u 1 2
Rp 1 2 1756
Cp 1 2 10.7p
Rs 1 N3 0.01
L1 N3 2 1.068u
.ends 5030_78438367010_1u
*******
.subckt 5030_78438367022_2.2u 1 2
Rp 1 2 3190
Cp 1 2 13.963p
Rs 1 N3 0.014
L1 N3 2 2.296u
.ends 5030_78438367022_2.2u
*******
.subckt 5030_78438367033_3.3u 1 2
Rp 1 2 4284
Cp 1 2 15.228p
Rs 1 N3 0.02
L1 N3 2 3.388u
.ends 5030_78438367033_3.3u
*******
.subckt 5030_78438367047_4.7u 1 2
Rp 1 2 5903
Cp 1 2 15.57p
Rs 1 N3 0.03
L1 N3 2 4.699u
.ends 5030_78438367047_4.7u
*******
.subckt 5030_78438367068_6.8u 1 2
Rp 1 2 7062
Cp 1 2 15.983p
Rs 1 N3 0.042
L1 N3 2 6.597u
.ends 5030_78438367068_6.8u
*******
.subckt 5030_78438367082_8.2u 1 2
Rp 1 2 6565
Cp 1 2 16.689p
Rs 1 N3 0.05
L1 N3 2 8.973u
.ends 5030_78438367082_8.2u
*******
.subckt 5030_78438367100_10u 1 2
Rp 1 2 7290
Cp 1 2 15.66p
Rs 1 N3 0.061
L1 N3 2 9.563u
.ends 5030_78438367100_10u
*******
.subckt 2010_784383430033_0.33u 1 2
Rp 1 2 1106.761952154
Cp 1 2 1.8829p
Rs 1 N3 0.04
L1 N3 2 0.32u
.ends 2010_784383430033_0.33u
*******
.subckt 2010_784383430047_0.47u 1 2
Rp 1 2 1457.590564128
Cp 1 2 1.9781p
Rs 1 N3 0.049
L1 N3 2 0.44u
.ends 2010_784383430047_0.47u
*******
.subckt 2010_784383430056_0.56u 1 2
Rp 1 2 2075.350512116
Cp 1 2 2.2551p
Rs 1 N3 0.056
L1 N3 2 0.5u
.ends 2010_784383430056_0.56u
*******
.subckt 2010_784383430068_0.68u 1 2
Rp 1 2 2110.665367845
Cp 1 2 2.1367p
Rs 1 N3 0.065
L1 N3 2 0.65u
.ends 2010_784383430068_0.68u
*******
.subckt 2010_784383430082_0.82u 1 2
Rp 1 2 2321.539322436
Cp 1 2 2.3941p
Rs 1 N3 0.071
L1 N3 2 0.76u
.ends 2010_784383430082_0.82u
*******
.subckt 2010_78438343010_1u 1 2
Rp 1 2 3024.486229762
Cp 1 2 2.6486p
Rs 1 N3 0.086
L1 N3 2 0.99u
.ends 2010_78438343010_1u
*******
.subckt 2010_78438343012_1.2u 1 2
Rp 1 2 3525.586090584
Cp 1 2 2.6299p
Rs 1 N3 0.114
L1 N3 2 1.07u
.ends 2010_78438343012_1.2u
*******
.subckt 2010_78438343015_1.5u 1 2
Rp 1 2 4272.400063088
Cp 1 2 2.4725p
Rs 1 N3 0.15
L1 N3 2 1.43u
.ends 2010_78438343015_1.5u
*******
.subckt 2010_78438343022_2.2u 1 2
Rp 1 2 5817.620850408
Cp 1 2 2.7082p
Rs 1 N3 0.225
L1 N3 2 1.92u
.ends 2010_78438343022_2.2u
*******
.subckt 4012_7843835400033_0.033u 1 2
Rp 1 2 157.464
Cp 1 2 1.69p
Rs 1 N3 0.0009
L1 N3 2 0.032211u
.ends 4012_7843835400033_0.033u
*******
.subckt 4012_7843835400068_0.068u 1 2
Rp 1 2 229.552
Cp 1 2 2.854p
Rs 1 N3 0.0017
L1 N3 2 0.063398u
.ends 4012_7843835400068_0.068u
*******
.subckt 2512HT_784383240033HT_0.33u 1 2
Rp 1 2 713.532
Cp 1 2 2.928p
Rs 1 N3 0.0232
L1 N3 2 0.286249u
.ends 2512HT_784383240033HT_0.33u
*******
.subckt 2512HT_784383240047HT_0.47u 1 2
Rp 1 2 1014
Cp 1 2 3.558p
Rs 1 N3 0.0301
L1 N3 2 0.412145u
.ends 2512HT_784383240047HT_0.47u
*******
.subckt 2512HT_784383240056HT_0.56u 1 2
Rp 1 2 1383
Cp 1 2 4.249p
Rs 1 N3 0.0383
L1 N3 2 0.567452u
.ends 2512HT_784383240056HT_0.56u
*******
.subckt 2512HT_78438324010HT_1u 1 2
Rp 1 2 2258
Cp 1 2 4.965p
Rs 1 N3 0.0534
L1 N3 2 1.015u
.ends 2512HT_78438324010HT_1u
*******
.subckt 2512HT_78438324012HT_1.2u 1 2
Rp 1 2 2590
Cp 1 2 4.76p
Rs 1 N3 0.0649
L1 N3 2 1.19u
.ends 2512HT_78438324012HT_1.2u
*******
.subckt 2512HT_78438324015HT_1.5u 1 2
Rp 1 2 3572
Cp 1 2 5.011p
Rs 1 N3 0.0887
L1 N3 2 1.606u
.ends 2512HT_78438324015HT_1.5u
*******
.subckt 2512HT_78438324022HT_2.2u 1 2
Rp 1 2 4359
Cp 1 2 4.441p
Rs 1 N3 0.1413
L1 N3 2 2.036u
.ends 2512HT_78438324022HT_2.2u
*******
.subckt 2512HT_78438324033HT_3.3u 1 2
Rp 1 2 5972
Cp 1 2 4.542p
Rs 1 N3 0.2388
L1 N3 2 3.179u
.ends 2512HT_78438324033HT_3.3u
*******
.subckt 2512HT_78438324047HT_4.7u 1 2
Rp 1 2 8027
Cp 1 2 5.136p
Rs 1 N3 0.3196
L1 N3 2 4.488u
.ends 2512HT_78438324047HT_4.7u
*******
.subckt 3015HT_784383350056HT_0.56u 1 2
Rp 1 2 1233
Cp 1 2 5.884p
Rs 1 N3 0.0193
L1 N3 2 0.494u
.ends 3015HT_784383350056HT_0.56u
*******
.subckt 3015HT_784383350068HT_0.68u 1 2
Rp 1 2 1632
Cp 1 2 6.41p
Rs 1 N3 0.0221
L1 N3 2 0.658u
.ends 3015HT_784383350068HT_0.68u
*******
.subckt 3015HT_78438335010HT_1u 1 2
Rp 1 2 2361
Cp 1 2 5.162p
Rs 1 N3 0.0462
L1 N3 2 0.925u
.ends 3015HT_78438335010HT_1u
*******
.subckt 3015HT_78438335022HT_2.2u 1 2
Rp 1 2 4091
Cp 1 2 7.078p
Rs 1 N3 0.0834
L1 N3 2 2.04u
.ends 3015HT_78438335022HT_2.2u
*******
.subckt 3015HT_78438335033HT_3.3u 1 2
Rp 1 2 6465
Cp 1 2 6.813p
Rs 1 N3 0.1156
L1 N3 2 3.01u
.ends 3015HT_78438335033HT_3.3u
*******
.subckt 3015HT_78438335047HT_4.7u 1 2
Rp 1 2 7862
Cp 1 2 7.621p
Rs 1 N3 0.1629
L1 N3 2 4.829u
.ends 3015HT_78438335047HT_4.7u
*******
.subckt 3015HT_78438335068HT_6.8u 1 2
Rp 1 2 9282
Cp 1 2 7.56p
Rs 1 N3 0.2701
L1 N3 2 6.915u
.ends 3015HT_78438335068HT_6.8u
*******
.subckt 3015HT_78438335100HT_10u 1 2
Rp 1 2 11568
Cp 1 2 8.042p
Rs 1 N3 0.4778
L1 N3 2 9.231u
.ends 3015HT_78438335100HT_10u
*******
.subckt 3020HT_784383360068HT_0.68u 1 2
Rp 1 2 1504
Cp 1 2 5.503p
Rs 1 N3 0.0244
L1 N3 2 0.636u
.ends 3020HT_784383360068HT_0.68u
*******
.subckt 3020HT_78438336010HT_1u 1 2
Rp 1 2 2123
Cp 1 2 5.792p
Rs 1 N3 0.0285
L1 N3 2 0.978u
.ends 3020HT_78438336010HT_1u
*******
.subckt 3020HT_78438336012HT_1.2u 1 2
Rp 1 2 2341
Cp 1 2 6.396p
Rs 1 N3 0.0326
L1 N3 2 1.119u
.ends 3020HT_78438336012HT_1.2u
*******
.subckt 3020HT_78438336015HT_1.5u 1 2
Rp 1 2 2851
Cp 1 2 6.152p
Rs 1 N3 0.0352
L1 N3 2 1.47u
.ends 3020HT_78438336015HT_1.5u
*******
.subckt 3020HT_78438336022HT_2.2u 1 2
Rp 1 2 4559
Cp 1 2 5.855p
Rs 1 N3 0.0569
L1 N3 2 1.952u
.ends 3020HT_78438336022HT_2.2u
*******
.subckt 3020HT_78438336033HT_3.3u 1 2
Rp 1 2 6126
Cp 1 2 6.307p
Rs 1 N3 0.0859
L1 N3 2 2.893u
.ends 3020HT_78438336033HT_3.3u
*******
.subckt 3020HT_78438336047HT_4.7u 1 2
Rp 1 2 7667
Cp 1 2 7.768p
Rs 1 N3 0.1306
L1 N3 2 4.215u
.ends 3020HT_78438336047HT_4.7u
*******
.subckt 3020HT_78438336068HT_6.8u 1 2
Rp 1 2 10703
Cp 1 2 8.277p
Rs 1 N3 0.1974
L1 N3 2 6.315u
.ends 3020HT_78438336068HT_6.8u
*******
.subckt 6030HT_784383770033HT_0.33u 1 2
Rp 1 2 666
Cp 1 2 8.985p
Rs 1 N3 0.0026
L1 N3 2 0.304u
.ends 6030HT_784383770033HT_0.33u
*******
.subckt 6030HT_784383770068HT_0.68u 1 2
Rp 1 2 1585
Cp 1 2 11.485p
Rs 1 N3 0.0048
L1 N3 2 0.728u
.ends 6030HT_784383770068HT_0.68u
*******
.subckt 6030HT_78438377010HT_1u 1 2
Rp 1 2 2159
Cp 1 2 11.644p
Rs 1 N3 0.006
L1 N3 2 0.981u
.ends 6030HT_78438377010HT_1u
*******
.subckt 6030HT_78438377022HT_2.2u 1 2
Rp 1 2 3944
Cp 1 2 15.465p
Rs 1 N3 0.0119
L1 N3 2 2.117u
.ends 6030HT_78438377022HT_2.2u
*******
.subckt 6030HT_78438377033HT_3.3u 1 2
Rp 1 2 5737
Cp 1 2 16.068p
Rs 1 N3 0.0177
L1 N3 2 3.253u
.ends 6030HT_78438377033HT_3.3u
*******
