**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  MLCCs - Multilayer Ceramic Chip Capacitors
* Matchcode:              WCAP-CSGP_6-3V
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/19/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0201_885012004011_10pF 1 2
Rser 1 3 0.5169
Lser 2 4 0.00000000022
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0201_885012004011_10pF
*******
.subckt 0201_885012004012_22pF 1 2
Rser 1 3 0.4505
Lser 2 4 0.000000000253
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0201_885012004012_22pF
*******
.subckt 0201_885012004013_33pF 1 2
Rser 1 3 0.2722
Lser 2 4 0.00000000022
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0201_885012004013_33pF
*******
.subckt 0201_885012004002_47pF 1 2
Rser 1 3 0.2226
Lser 2 4 0.0000000002
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0201_885012004002_47pF
*******
.subckt 0201_885012204001_100pF 1 2
Rser 1 3 0.8951
Lser 2 4 0.00000000017
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0201_885012204001_100pF
*******
.subckt 0201_885012004014_100pF 1 2
Rser 1 3 0.1789
Lser 2 4 0.0000000002
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0201_885012004014_100pF
*******
.subckt 0201_885012204002_680pF 1 2
Rser 1 3 0.3189
Lser 2 4 0.00000000022
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0201_885012204002_680pF
*******
.subckt 0201_885012204003_1nF 1 2
Rser 1 3 0.2506
Lser 2 4 0.00000000021
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0201_885012204003_1nF
*******
.subckt 0402_885012005049_1pF 1 2
Rser 1 3 0.372412566115
Lser 2 4 3.42487064E-10
C1 3 4 0.000000000001
Rpar 3 4 10000000000
.ends 0402_885012005049_1pF
*******
.subckt 0402_885012005050_1.5pF 1 2
Rser 1 3 1.6
Lser 2 4 0.00000000034
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0402_885012005050_1.5pF
*******
.subckt 0402_885012005051_2.2pF 1 2
Rser 1 3 0.373107051593
Lser 2 4 3.52926651E-10
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0402_885012005051_2.2pF
*******
.subckt 0402_885012005052_3.3pF 1 2
Rser 1 3 0.7
Lser 2 4 0.0000000004
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0402_885012005052_3.3pF
*******
.subckt 0402_885012005053_4.7pF 1 2
Rser 1 3 0.443688812845
Lser 2 4 4.55408482E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0402_885012005053_4.7pF
*******
.subckt 0402_885012005054_6.8pF 1 2
Rser 1 3 0.397780736645
Lser 2 4 4.18761945E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0402_885012005054_6.8pF
*******
.subckt 0402_885012005055_10pF 1 2
Rser 1 3 0.367986500147
Lser 2 4 4.54592782E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005055_10pF
*******
.subckt 0402_885012005056_15pF 1 2
Rser 1 3 0.289002377009
Lser 2 4 4.35524241E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0402_885012005056_15pF
*******
.subckt 0402_885012005057_22pF 1 2
Rser 1 3 0.1946461244
Lser 2 4 4.43759844E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0402_885012005057_22pF
*******
.subckt 0402_885012005058_33pF 1 2
Rser 1 3 0.125165063018
Lser 2 4 4.11479308E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005058_33pF
*******
.subckt 0402_885012005059_47pF 1 2
Rser 1 3 0.136483462277
Lser 2 4 4.44322285E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005059_47pF
*******
.subckt 0402_885012005060_68pF 1 2
Rser 1 3 0.101411214779
Lser 2 4 4.24748886E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005060_68pF
*******
.subckt 0402_885012005061_100pF 1 2
Rser 1 3 0.0708016190464
Lser 2 4 3.72654022E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005061_100pF
*******
.subckt 0402_885012005062_150pF 1 2
Rser 1 3 0.043551770519
Lser 2 4 3.72165147E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012005062_150pF
*******
.subckt 0402_885012005063_220pF 1 2
Rser 1 3 0.0328677075671
Lser 2 4 3.55619232E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012005063_220pF
*******
.subckt 0402_885012005067_1nF 1 2
Rser 1 3 0.127
Lser 2 4 1.020979922E-09
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012005067_1nF
*******
.subckt 0402_885012205055_100pF 1 2
Rser 1 3 0.81826
Lser 2 4 0.00000000027428
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012205055_100pF
*******
.subckt 0402_885012205056_150pF 1 2
Rser 1 3 0.632711426036
Lser 2 4 1.20280732E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0402_885012205056_150pF
*******
.subckt 0402_885012205057_220pF 1 2
Rser 1 3 0.578964014005
Lser 2 4 1.69232145E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0402_885012205057_220pF
*******
.subckt 0402_885012205058_330pF 1 2
Rser 1 3 0.503553103715
Lser 2 4 1.67673778E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0402_885012205058_330pF
*******
.subckt 0402_885012205059_470pF 1 2
Rser 1 3 0.341891187733
Lser 2 4 1.53352894E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0402_885012205059_470pF
*******
.subckt 0402_885012205060_680pF 1 2
Rser 1 3 0.291776877274
Lser 2 4 1.90727531E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0402_885012205060_680pF
*******
.subckt 0402_885012205061_1nF 1 2
Rser 1 3 0.16682
Lser 2 4 0.00000000027542
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205061_1nF
*******
.subckt 0402_885012205062_1.5nF 1 2
Rser 1 3 0.318149132739
Lser 2 4 2.00030416E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0402_885012205062_1.5nF
*******
.subckt 0402_885012205063_2.2nF 1 2
Rser 1 3 0.167940534432
Lser 2 4 1.9652905E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0402_885012205063_2.2nF
*******
.subckt 0402_885012205064_3.3nF 1 2
Rser 1 3 0.128032535119
Lser 2 4 2.21229721E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0402_885012205064_3.3nF
*******
.subckt 0402_885012205065_4.7nF 1 2
Rser 1 3 0.12665496656
Lser 2 4 2.40553052E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205065_4.7nF
*******
.subckt 0402_885012205066_6.8nF 1 2
Rser 1 3 0.103789689499
Lser 2 4 1.90645336E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0402_885012205066_6.8nF
*******
.subckt 0402_885012205067_10nF 1 2
Rser 1 3 0.110942181295
Lser 2 4 1.63617133E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0402_885012205067_10nF
*******
.subckt 0402_885012205086_100nF 1 2
Rser 1 3 0.07
Lser 2 4 0.00000000055
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0402_885012205086_100nF
*******
.subckt 0402_885012205092_100nF 1 2
Rser 1 3 0.033
Lser 2 4 0.0000000006
C1 3 4 0.0000001
Rpar 3 4 500000000
.ends 0402_885012205092_100nF
*******
.subckt 0603_885012006048_3.3pF 1 2
Rser 1 3 0.351777802818
Lser 2 4 4.93521689E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0603_885012006048_3.3pF
*******
.subckt 0603_885012006049_4.7pF 1 2
Rser 1 3 0.314951809581
Lser 2 4 4.34213899E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0603_885012006049_4.7pF
*******
.subckt 0603_885012006050_6.8pF 1 2
Rser 1 3 0.53
Lser 2 4 0.00000000049
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0603_885012006050_6.8pF
*******
.subckt 0603_885012006051_10pF 1 2
Rser 1 3 0.423568844547
Lser 2 4 6.08699424E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006051_10pF
*******
.subckt 0603_885012006052_15pF 1 2
Rser 1 3 0.396040749585
Lser 2 4 6.08298711E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006052_15pF
*******
.subckt 0603_885012006053_22pF 1 2
Rser 1 3 0.388744823765
Lser 2 4 6.9588017E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006053_22pF
*******
.subckt 0603_885012006054_33pF 1 2
Rser 1 3 0.321193198235
Lser 2 4 7.31689517E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006054_33pF
*******
.subckt 0603_885012006055_47pF 1 2
Rser 1 3 0.290935011258
Lser 2 4 4.02698987E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006055_47pF
*******
.subckt 0603_885012006056_68pF 1 2
Rser 1 3 0.190199312239
Lser 2 4 6.75111985E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006056_68pF
*******
.subckt 0603_885012006057_100pF 1 2
Rser 1 3 0.155626039874
Lser 2 4 4.37579661E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006057_100pF
*******
.subckt 0603_885012006058_150pF 1 2
Rser 1 3 0.117171082106
Lser 2 4 5.86950362E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006058_150pF
*******
.subckt 0603_885012006059_220pF 1 2
Rser 1 3 0.120673949599
Lser 2 4 6.11171216E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012006059_220pF
*******
.subckt 0603_885012006060_330pF 1 2
Rser 1 3 0.0984499950001
Lser 2 4 5.75039775E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006060_330pF
*******
.subckt 0603_885012006061_470pF 1 2
Rser 1 3 0.0701665420081
Lser 2 4 5.55279727E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006061_470pF
*******
.subckt 0603_885012006062_680pF 1 2
Rser 1 3 0.058780576404
Lser 2 4 5.07120306E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006062_680pF
*******
.subckt 0603_885012006063_1nF 1 2
Rser 1 3 0.040317449025
Lser 2 4 4.45418718E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006063_1nF
*******
.subckt 0603_885012006094_100pF 1 2
Rser 1 3 0.149672201927
Lser 2 4 1.208801635E-09
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006094_100pF
*******
.subckt 0603_885012006096_150pF 1 2
Rser 1 3 0.119
Lser 2 4 0.00000000118
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006096_150pF
*******
.subckt 0603_885012006097_1nF 1 2
Rser 1 3 0.0539689392343
Lser 2 4 1.060354109E-09
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006097_1nF
*******
.subckt 0603_885012206077_100pF 1 2
Rser 1 3 0.85996
Lser 2 4 0.00000000023099
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206077_100pF
*******
.subckt 0603_885012206078_150pF 1 2
Rser 1 3 0.6711
Lser 2 4 0.00000000028059
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012206078_150pF
*******
.subckt 0603_885012206079_220pF 1 2
Rser 1 3 0.58208
Lser 2 4 0.00000000030164
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0603_885012206079_220pF
*******
.subckt 0603_885012206080_330pF 1 2
Rser 1 3 0.43473
Lser 2 4 0.00000000032084
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206080_330pF
*******
.subckt 0603_885012206081_470pF 1 2
Rser 1 3 0.34619
Lser 2 4 0.00000000032738
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206081_470pF
*******
.subckt 0603_885012206082_680pF 1 2
Rser 1 3 0.303992916785
Lser 2 4 3.80425244E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206082_680pF
*******
.subckt 0603_885012206083_1nF 1 2
Rser 1 3 0.25783718447
Lser 2 4 4.104475E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206083_1nF
*******
.subckt 0603_885012206084_1.5nF 1 2
Rser 1 3 0.180999474852
Lser 2 4 3.54773595E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206084_1.5nF
*******
.subckt 0603_885012206085_2.2nF 1 2
Rser 1 3 0.139424404216
Lser 2 4 3.27512531E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0603_885012206085_2.2nF
*******
.subckt 0603_885012206086_3.3nF 1 2
Rser 1 3 0.105745225203
Lser 2 4 3.39462116E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206086_3.3nF
*******
.subckt 0603_885012206087_4.7nF 1 2
Rser 1 3 0.0821607581427
Lser 2 4 2.83989011E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206087_4.7nF
*******
.subckt 0603_885012206088_6.8nF 1 2
Rser 1 3 0.0838686105847
Lser 2 4 4.16447222E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206088_6.8nF
*******
.subckt 0603_885012206089_10nF 1 2
Rser 1 3 0.0358532866879
Lser 2 4 3.4059544E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206089_10nF
*******
.subckt 0603_885012206090_15nF 1 2
Rser 1 3 0.0485012368007
Lser 2 4 3.32575255E-10
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0603_885012206090_15nF
*******
.subckt 0603_885012206091_22nF 1 2
Rser 1 3 0.00971971773084
Lser 2 4 3.00225265E-10
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0603_885012206091_22nF
*******
.subckt 0603_885012206092_33nF 1 2
Rser 1 3 0.02322
Lser 2 4 0.00000000030071
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0603_885012206092_33nF
*******
.subckt 0603_885012206093_47nF 1 2
Rser 1 3 0.02723
Lser 2 4 0.00000000027891
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0603_885012206093_47nF
*******
.subckt 0603_885012206094_68nF 1 2
Rser 1 3 0.01852
Lser 2 4 0.00000000023609
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0603_885012206094_68nF
*******
.subckt 0603_885012206095_100nF 1 2
Rser 1 3 0.0157659152881
Lser 2 4 3.10171966E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206095_100nF
*******
.subckt 0603_885012206121_330nF 1 2
Rser 1 3 0.0116331902783
Lser 2 4 2.98906197E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0603_885012206121_330nF
*******
.subckt 0603_885012206125_220nF 1 2
Rser 1 3 0.017
Lser 2 4 0.000000001
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0603_885012206125_220nF
*******
.subckt 0603_885012206126_1uF 1 2
Rser 1 3 0.0115
Lser 2 4 0.0000000008
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 0603_885012206126_1uF
*******
.subckt 0603_885012206083R_1nF 1 2
Rser 1 3 0.25783718447
Lser 2 4 4.104475E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206083R_1nF
*******
.subckt 0603_885012206089R_10nF 1 2
Rser 1 3 0.0358532866879
Lser 2 4 3.4059544E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206089R_10nF
*******
.subckt 0603_885012206095R_100nF 1 2
Rser 1 3 0.0157659152881
Lser 2 4 3.10171966E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0603_885012206095R_100nF
*******
.subckt 0603_885012006095_22pF 1 2
Rser 1 3 0.022
Lser 2 4 0.0000000011
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0603_885012006095_22pF
*******
.subckt 0805_885012007046_1.5pF 1 2
Rser 1 3 0.498754904967
Lser 2 4 4.46307458E-10
C1 3 4 0.0000000000015
Rpar 3 4 10000000000
.ends 0805_885012007046_1.5pF
*******
.subckt 0805_885012007047_2.2pF 1 2
Rser 1 3 0.464027184378
Lser 2 4 4.17958974E-10
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0805_885012007047_2.2pF
*******
.subckt 0805_885012007048_3.3pF 1 2
Rser 1 3 0.476983731701
Lser 2 4 4.57833988E-10
C1 3 4 0.0000000000033
Rpar 3 4 10000000000
.ends 0805_885012007048_3.3pF
*******
.subckt 0805_885012007049_4.7pF 1 2
Rser 1 3 0.497100489266
Lser 2 4 4.97943432E-10
C1 3 4 0.0000000000047
Rpar 3 4 10000000000
.ends 0805_885012007049_4.7pF
*******
.subckt 0805_885012007050_6.8pF 1 2
Rser 1 3 0.437292047874
Lser 2 4 5.43803179E-10
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 0805_885012007050_6.8pF
*******
.subckt 0805_885012007051_10pF 1 2
Rser 1 3 0.5317
Lser 2 4 0.00000000045
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0805_885012007051_10pF
*******
.subckt 0805_885012007052_15pF 1 2
Rser 1 3 0.351715326777
Lser 2 4 5.44262413E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007052_15pF
*******
.subckt 0805_885012007053_22pF 1 2
Rser 1 3 0.320807516938
Lser 2 4 5.98353392E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 0805_885012007053_22pF
*******
.subckt 0805_885012007054_33pF 1 2
Rser 1 3 0.251170142371
Lser 2 4 5.67157711E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007054_33pF
*******
.subckt 0805_885012007055_47pF 1 2
Rser 1 3 0.216515950035
Lser 2 4 5.20835554E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885012007055_47pF
*******
.subckt 0805_885012007056_68pF 1 2
Rser 1 3 0.173987704202
Lser 2 4 4.36318354E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0805_885012007056_68pF
*******
.subckt 0805_885012007057_100pF 1 2
Rser 1 3 0.112239658687
Lser 2 4 3.23857063E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007057_100pF
*******
.subckt 0805_885012007058_150pF 1 2
Rser 1 3 0.125944924272
Lser 2 4 4.46129224E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007058_150pF
*******
.subckt 0805_885012007059_220pF 1 2
Rser 1 3 0.079249932999
Lser 2 4 3.92377309E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012007059_220pF
*******
.subckt 0805_885012007060_330pF 1 2
Rser 1 3 0.0873115639161
Lser 2 4 4.48869509E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007060_330pF
*******
.subckt 0805_885012007061_470pF 1 2
Rser 1 3 0.0447460793708
Lser 2 4 5.13925095E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007061_470pF
*******
.subckt 0805_885012007062_680pF 1 2
Rser 1 3 0.0641329981739
Lser 2 4 4.25300517E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012007062_680pF
*******
.subckt 0805_885012007063_1nF 1 2
Rser 1 3 0.0594421507531
Lser 2 4 4.12205624E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007063_1nF
*******
.subckt 0805_885012007064_1.5nF 1 2
Rser 1 3 0.0542761813318
Lser 2 4 4.44523189E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012007064_1.5nF
*******
.subckt 0805_885012007065_2.2nF 1 2
Rser 1 3 0.0452125293188
Lser 2 4 3.18286842E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012007065_2.2nF
*******
.subckt 0805_885012007066_3.3nF 1 2
Rser 1 3 0.0386718470366
Lser 2 4 4.52637868E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012007066_3.3nF
*******
.subckt 0805_885012007067_4.7nF 1 2
Rser 1 3 0.0321239026517
Lser 2 4 3.90170133E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012007067_4.7nF
*******
.subckt 0805_885012007105_470pF 1 2
Rser 1 3 0.07
Lser 2 4 0.0000000011
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007105_470pF
*******
.subckt 0805_885012007106_2.2nF 1 2
Rser 1 3 0.0409413211003
Lser 2 4 1.060592085E-09
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012007106_2.2nF
*******
.subckt 0805_885012007107_330pF 1 2
Rser 1 3 0.083
Lser 2 4 0.00000000106
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007107_330pF
*******
.subckt 0805_885012207080_100pF 1 2
Rser 1 3 0.88248
Lser 2 4 0.00000000026383
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207080_100pF
*******
.subckt 0805_885012207081_150pF 1 2
Rser 1 3 0.74128
Lser 2 4 0.00000000030962
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012207081_150pF
*******
.subckt 0805_885012207082_220pF 1 2
Rser 1 3 0.48326
Lser 2 4 0.00000000027382
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 0805_885012207082_220pF
*******
.subckt 0805_885012207083_330pF 1 2
Rser 1 3 0.40314
Lser 2 4 0.00000000028019
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012207083_330pF
*******
.subckt 0805_885012207084_470pF 1 2
Rser 1 3 0.29801
Lser 2 4 0.00000000032037
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207084_470pF
*******
.subckt 0805_885012207085_680pF 1 2
Rser 1 3 0.24191
Lser 2 4 0.00000000035763
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012207085_680pF
*******
.subckt 0805_885012207086_1nF 1 2
Rser 1 3 0.16468
Lser 2 4 0.00000000030011
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207086_1nF
*******
.subckt 0805_885012207087_1.5nF 1 2
Rser 1 3 0.14696
Lser 2 4 0.00000000040084
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207087_1.5nF
*******
.subckt 0805_885012207088_2.2nF 1 2
Rser 1 3 0.11179
Lser 2 4 0.00000000038067
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 0805_885012207088_2.2nF
*******
.subckt 0805_885012207089_3.3nF 1 2
Rser 1 3 0.08492
Lser 2 4 0.0000000003695
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207089_3.3nF
*******
.subckt 0805_885012207090_4.7nF 1 2
Rser 1 3 0.05225
Lser 2 4 0.00000000025076
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012207090_4.7nF
*******
.subckt 0805_885012207091_6.8nF 1 2
Rser 1 3 0.06481
Lser 2 4 0.00000000034495
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0805_885012207091_6.8nF
*******
.subckt 0805_885012207092_10nF 1 2
Rser 1 3 0.06275
Lser 2 4 0.00000000031024
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207092_10nF
*******
.subckt 0805_885012207093_15nF 1 2
Rser 1 3 0.04594
Lser 2 4 0.00000000031216
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 0805_885012207093_15nF
*******
.subckt 0805_885012207094_22nF 1 2
Rser 1 3 0.04966
Lser 2 4 0.00000000031956
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 0805_885012207094_22nF
*******
.subckt 0805_885012207095_33nF 1 2
Rser 1 3 0.0344549798517
Lser 2 4 0.00000000043
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 0805_885012207095_33nF
*******
.subckt 0805_885012207096_47nF 1 2
Rser 1 3 0.0256748827303
Lser 2 4 0.00000000038
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 0805_885012207096_47nF
*******
.subckt 0805_885012207097_68nF 1 2
Rser 1 3 0.0207501013107
Lser 2 4 0.00000000038
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 0805_885012207097_68nF
*******
.subckt 0805_885012207098_100nF 1 2
Rser 1 3 0.0175748078756
Lser 2 4 0.0000000004
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207098_100nF
*******
.subckt 0805_885012207099_150nF 1 2
Rser 1 3 0.0142447362747
Lser 2 4 0.00000000045
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 0805_885012207099_150nF
*******
.subckt 0805_885012207100_220nF 1 2
Rser 1 3 0.0120359560176
Lser 2 4 0.00000000044
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 0805_885012207100_220nF
*******
.subckt 0805_885012207101_330nF 1 2
Rser 1 3 0.0111899844274
Lser 2 4 0.00000000048
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 0805_885012207101_330nF
*******
.subckt 0805_885012207102_470nF 1 2
Rser 1 3 0.00874819634126
Lser 2 4 0.000000000465
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 0805_885012207102_470nF
*******
.subckt 0805_885012207103_1uF 1 2
Rser 1 3 0.0053065272233
Lser 2 4 2.83466289E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0805_885012207103_1uF
*******
.subckt 0805_885012207098R_100nF 1 2
Rser 1 3 0.0175748078756
Lser 2 4 0.0000000004
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 0805_885012207098R_100nF
*******
.subckt 0805_885012207103R_1uF 1 2
Rser 1 3 0.0053065272233
Lser 2 4 2.83466289E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 0805_885012207103R_1uF
*******
.subckt 1206_885012008036_6.8pF 1 2
Rser 1 3 0.37597
Lser 2 4 0.00000000066
C1 3 4 0.0000000000068
Rpar 3 4 10000000000
.ends 1206_885012008036_6.8pF
*******
.subckt 1206_885012008037_10pF 1 2
Rser 1 3 0.247786722229
Lser 2 4 5.75498755E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1206_885012008037_10pF
*******
.subckt 1206_885012008038_15pF 1 2
Rser 1 3 0.203981995296
Lser 2 4 5.79093876E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 1206_885012008038_15pF
*******
.subckt 1206_885012008039_22pF 1 2
Rser 1 3 0.160102464353
Lser 2 4 5.19970978E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1206_885012008039_22pF
*******
.subckt 1206_885012008040_33pF 1 2
Rser 1 3 0.211299340525
Lser 2 4 5.80360065E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 1206_885012008040_33pF
*******
.subckt 1206_885012008041_47pF 1 2
Rser 1 3 0.208069659743
Lser 2 4 5.31192815E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885012008041_47pF
*******
.subckt 1206_885012008042_68pF 1 2
Rser 1 3 0.207112222887
Lser 2 4 5.32291452E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 1206_885012008042_68pF
*******
.subckt 1206_885012008043_100pF 1 2
Rser 1 3 0.120593750684
Lser 2 4 4.75662979E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008043_100pF
*******
.subckt 1206_885012008044_150pF 1 2
Rser 1 3 0.116934479556
Lser 2 4 4.79036564E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012008044_150pF
*******
.subckt 1206_885012008045_220pF 1 2
Rser 1 3 0.10386657318
Lser 2 4 4.26569823E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012008045_220pF
*******
.subckt 1206_885012008046_330pF 1 2
Rser 1 3 0.0889473100116
Lser 2 4 3.86799658E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012008046_330pF
*******
.subckt 1206_885012008047_470pF 1 2
Rser 1 3 0.112293156509
Lser 2 4 4.49592146E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012008047_470pF
*******
.subckt 1206_885012008048_680pF 1 2
Rser 1 3 0.0885483556492
Lser 2 4 4.83404689E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012008048_680pF
*******
.subckt 1206_885012008049_1nF 1 2
Rser 1 3 0.0678258865879
Lser 2 4 4.38251746E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012008049_1nF
*******
.subckt 1206_885012008050_1.5nF 1 2
Rser 1 3 0.066
Lser 2 4 0.00000000118
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012008050_1.5nF
*******
.subckt 1206_885012008051_2.2nF 1 2
Rser 1 3 0.0481287677862
Lser 2 4 4.23334149E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012008051_2.2nF
*******
.subckt 1206_885012008052_3.3nF 1 2
Rser 1 3 0.048551433153
Lser 2 4 3.89367659E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012008052_3.3nF
*******
.subckt 1206_885012008053_4.7nF 1 2
Rser 1 3 0.0373751695173
Lser 2 4 3.96656883E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012008053_4.7nF
*******
.subckt 1206_885012008054_6.8nF 1 2
Rser 1 3 0.0328755784645
Lser 2 4 4.18880071E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008054_6.8nF
*******
.subckt 1206_885012008055_10nF 1 2
Rser 1 3 0.0308699044735
Lser 2 4 4.5821325E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008055_10nF
*******
.subckt 1206_885012008082_3.3nF 1 2
Rser 1 3 0.0433164856935
Lser 2 4 1.256573444E-09
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012008082_3.3nF
*******
.subckt 1206_885012108022_10uF 1 2
Rser 1 3 0.00342327531378
Lser 2 4 0.000000000799
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1206_885012108022_10uF
*******
.subckt 1206_885012208070_150pF 1 2
Rser 1 3 0.71274
Lser 2 4 0.00000000032053
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012208070_150pF
*******
.subckt 1206_885012208071_220pF 1 2
Rser 1 3 0.50529569726
Lser 2 4 2.96273344E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1206_885012208071_220pF
*******
.subckt 1206_885012208072_330pF 1 2
Rser 1 3 0.43202
Lser 2 4 0.00000000057877
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012208072_330pF
*******
.subckt 1206_885012208073_470pF 1 2
Rser 1 3 0.34146
Lser 2 4 0.00000000040636
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208073_470pF
*******
.subckt 1206_885012208074_680pF 1 2
Rser 1 3 0.34068
Lser 2 4 0.00000000050397
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012208074_680pF
*******
.subckt 1206_885012208075_1nF 1 2
Rser 1 3 0.22519
Lser 2 4 0.00000000041699
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208075_1nF
*******
.subckt 1206_885012208076_1.5nF 1 2
Rser 1 3 0.18074
Lser 2 4 0.00000000040041
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012208076_1.5nF
*******
.subckt 1206_885012208077_2.2nF 1 2
Rser 1 3 0.13842
Lser 2 4 0.00000000039067
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1206_885012208077_2.2nF
*******
.subckt 1206_885012208078_3.3nF 1 2
Rser 1 3 0.13733
Lser 2 4 0.00000000045693
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012208078_3.3nF
*******
.subckt 1206_885012208079_4.7nF 1 2
Rser 1 3 0.09403
Lser 2 4 0.00000000040583
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208079_4.7nF
*******
.subckt 1206_885012208080_6.8nF 1 2
Rser 1 3 0.08271
Lser 2 4 0.00000000048076
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012208080_6.8nF
*******
.subckt 1206_885012208081_10nF 1 2
Rser 1 3 0.07548
Lser 2 4 0.00000000050044
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208081_10nF
*******
.subckt 1206_885012208082_15nF 1 2
Rser 1 3 0.06346
Lser 2 4 0.00000000050869
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1206_885012208082_15nF
*******
.subckt 1206_885012208083_22nF 1 2
Rser 1 3 0.05996
Lser 2 4 0.00000000050024
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1206_885012208083_22nF
*******
.subckt 1206_885012208084_33nF 1 2
Rser 1 3 0.07214
Lser 2 4 0.00000000048096
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1206_885012208084_33nF
*******
.subckt 1206_885012208085_47nF 1 2
Rser 1 3 0.05144
Lser 2 4 0.00000000044024
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1206_885012208085_47nF
*******
.subckt 1206_885012208086_68nF 1 2
Rser 1 3 0.03887
Lser 2 4 0.00000000042372
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 1206_885012208086_68nF
*******
.subckt 1206_885012208087_100nF 1 2
Rser 1 3 0.02357
Lser 2 4 0.00000000059109
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1206_885012208087_100nF
*******
.subckt 1206_885012208088_150nF 1 2
Rser 1 3 0.01669
Lser 2 4 0.00000000057596
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1206_885012208088_150nF
*******
.subckt 1206_885012208089_220nF 1 2
Rser 1 3 0.01154
Lser 2 4 0.0000000005471
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1206_885012208089_220nF
*******
.subckt 1206_885012208090_330nF 1 2
Rser 1 3 0.01154
Lser 2 4 0.00000000068941
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1206_885012208090_330nF
*******
.subckt 1206_885012208091_470nF 1 2
Rser 1 3 0.01065
Lser 2 4 0.00000000073215
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1206_885012208091_470nF
*******
.subckt 1206_885012208092_680nF 1 2
Rser 1 3 0.00829
Lser 2 4 0.00000000068878
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1206_885012208092_680nF
*******
.subckt 1206_885012208093_1uF 1 2
Rser 1 3 0.00556
Lser 2 4 0.00000000059996
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1206_885012208093_1uF
*******
.subckt 1206_885012208094_4.7uF 1 2
Rser 1 3 0.00352
Lser 2 4 0.00000000057332
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1206_885012208094_4.7uF
*******
.subckt 1210_885012009007_22pF 1 2
Rser 1 3 0.374121714519
Lser 2 4 2.35270135E-10
C1 3 4 0.000000000022
Rpar 3 4 10000000000
.ends 1210_885012009007_22pF
*******
.subckt 1210_885012009008_33pF 1 2
Rser 1 3 0.242364797292
Lser 2 4 2.04183536E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 1210_885012009008_33pF
*******
.subckt 1210_885012009009_47pF 1 2
Rser 1 3 0.210290362797
Lser 2 4 2.1842961E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1210_885012009009_47pF
*******
.subckt 1210_885012009010_68pF 1 2
Rser 1 3 0.147762447298
Lser 2 4 1.90656729E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 1210_885012009010_68pF
*******
.subckt 1210_885012009011_100pF 1 2
Rser 1 3 0.129347366442
Lser 2 4 2.02608781E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1210_885012009011_100pF
*******
.subckt 1210_885012009012_150pF 1 2
Rser 1 3 0.130052835884
Lser 2 4 2.16784494E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1210_885012009012_150pF
*******
.subckt 1210_885012009013_220pF 1 2
Rser 1 3 0.0421105658392
Lser 2 4 2.03486371E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1210_885012009013_220pF
*******
.subckt 1210_885012009014_330pF 1 2
Rser 1 3 0.0366680474844
Lser 2 4 2.12935248E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1210_885012009014_330pF
*******
.subckt 1210_885012009015_470pF 1 2
Rser 1 3 0.041753756573
Lser 2 4 3.51053092E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1210_885012009015_470pF
*******
.subckt 1210_885012009016_680pF 1 2
Rser 1 3 0.0310627645209
Lser 2 4 2.06977272E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1210_885012009016_680pF
*******
.subckt 1210_885012009017_1nF 1 2
Rser 1 3 0.0212060307253
Lser 2 4 2.0371621E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885012009017_1nF
*******
.subckt 1210_885012009018_1.5nF 1 2
Rser 1 3 0.0312392079081
Lser 2 4 2.87207915E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1210_885012009018_1.5nF
*******
.subckt 1210_885012009019_2.2nF 1 2
Rser 1 3 0.0215418747712
Lser 2 4 2.06777607E-10
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1210_885012009019_2.2nF
*******
.subckt 1210_885012009020_3.3nF 1 2
Rser 1 3 0.0267047192368
Lser 2 4 2.05676794E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1210_885012009020_3.3nF
*******
.subckt 1210_885012009021_4.7nF 1 2
Rser 1 3 0.0311921178887
Lser 2 4 2.6092549E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1210_885012009021_4.7nF
*******
.subckt 1210_885012009022_6.8nF 1 2
Rser 1 3 0.0328474651911
Lser 2 4 1.68986675E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1210_885012009022_6.8nF
*******
.subckt 1210_885012009023_10nF 1 2
Rser 1 3 0.0123831418384
Lser 2 4 1.88456734E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1210_885012009023_10nF
*******
.subckt 1210_885012009024_15nF 1 2
Rser 1 3 0.0151582048451
Lser 2 4 2.71190675E-10
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1210_885012009024_15nF
*******
.subckt 1210_885012209029_1nF 1 2
Rser 1 3 0.24578
Lser 2 4 0.00000000010314
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1210_885012209029_1nF
*******
.subckt 1210_885012209030_1.5nF 1 2
Rser 1 3 0.21363
Lser 2 4 0.00000000011258
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1210_885012209030_1.5nF
*******
.subckt 1210_885012209031_2.2nF 1 2
Rser 1 3 0.17328
Lser 2 4 0.00000000013551
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1210_885012209031_2.2nF
*******
.subckt 1210_885012209032_3.3nF 1 2
Rser 1 3 0.10148
Lser 2 4 0.000000000079128
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1210_885012209032_3.3nF
*******
.subckt 1210_885012209033_4.7nF 1 2
Rser 1 3 0.12905
Lser 2 4 0.00000000012069
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1210_885012209033_4.7nF
*******
.subckt 1210_885012209034_6.8nF 1 2
Rser 1 3 0.05767
Lser 2 4 0.0000000001329
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1210_885012209034_6.8nF
*******
.subckt 1210_885012209035_10nF 1 2
Rser 1 3 0.07029
Lser 2 4 0.00000000063234
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1210_885012209035_10nF
*******
.subckt 1210_885012209036_15nF 1 2
Rser 1 3 0.04823
Lser 2 4 0.00000000065476
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1210_885012209036_15nF
*******
.subckt 1210_885012209037_22nF 1 2
Rser 1 3 0.0318
Lser 2 4 0.0000000005907
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1210_885012209037_22nF
*******
.subckt 1210_885012209038_33nF 1 2
Rser 1 3 0.02862
Lser 2 4 0.00000000012573
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1210_885012209038_33nF
*******
.subckt 1210_885012209039_47nF 1 2
Rser 1 3 0.01636
Lser 2 4 0.00000000055283
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1210_885012209039_47nF
*******
.subckt 1210_885012209040_68nF 1 2
Rser 1 3 0.02967
Lser 2 4 0.00000000066933
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 1210_885012209040_68nF
*******
.subckt 1210_885012209041_100nF 1 2
Rser 1 3 0.0232640980559
Lser 2 4 5.50483551E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1210_885012209041_100nF
*******
.subckt 1210_885012209042_150nF 1 2
Rser 1 3 0.0151905172405
Lser 2 4 5.27589443E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1210_885012209042_150nF
*******
.subckt 1210_885012209043_220nF 1 2
Rser 1 3 0.0127857665848
Lser 2 4 5.1481312E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1210_885012209043_220nF
*******
.subckt 1210_885012209044_330nF 1 2
Rser 1 3 0.00839371610696
Lser 2 4 5.53587415E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1210_885012209044_330nF
*******
.subckt 1210_885012209045_470nF 1 2
Rser 1 3 0.00675106116736
Lser 2 4 5.53881923E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1210_885012209045_470nF
*******
.subckt 1210_885012209046_680nF 1 2
Rser 1 3 0.00595213609047
Lser 2 4 5.69870142E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1210_885012209046_680nF
*******
.subckt 1210_885012209047_1uF 1 2
Rser 1 3 0.0444403254894
Lser 2 4 7.99001148E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209047_1uF
*******
.subckt 1210_885012209048_4.7uF 1 2
Rser 1 3 0.00278836774782
Lser 2 4 2.60340728E-10
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 1210_885012209048_4.7uF
*******
.subckt 1210_885012209073_10uF 1 2
Rser 1 3 0.00803494307495
Lser 2 4 4.01881911E-10
C1 3 4 0.00001
Rpar 3 4 5000000
.ends 1210_885012209073_10uF
*******
.subckt 1210_885012209047R_1uF 1 2
Rser 1 3 0.0444403254894
Lser 2 4 7.99001148E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1210_885012209047R_1uF
*******
.subckt 1812_885012010005_100pF 1 2
Rser 1 3 0.12355169432
Lser 2 4 3.51203653E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1812_885012010005_100pF
*******
.subckt 1812_885012010006_220pF 1 2
Rser 1 3 0.0878558292315
Lser 2 4 3.98601571E-10
C1 3 4 0.00000000022
Rpar 3 4 10000000000
.ends 1812_885012010006_220pF
*******
.subckt 1812_885012010007_470pF 1 2
Rser 1 3 0.0486179980779
Lser 2 4 3.42708418E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1812_885012010007_470pF
*******
.subckt 1812_885012010008_1nF 1 2
Rser 1 3 0.054974361057
Lser 2 4 3.20553197E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_885012010008_1nF
*******
.subckt 1812_885012010009_1.5nF 1 2
Rser 1 3 0.0235411944876
Lser 2 4 3.17035352E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1812_885012010009_1.5nF
*******
.subckt 1812_885012010010_3.3nF 1 2
Rser 1 3 0.0199944630408
Lser 2 4 3.02916593E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1812_885012010010_3.3nF
*******
.subckt 1812_885012010011_4.7nF 1 2
Rser 1 3 0.0944854934425
Lser 2 4 4.17148603E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1812_885012010011_4.7nF
*******
.subckt 1812_885012010012_6.8nF 1 2
Rser 1 3 0.0862794087323
Lser 2 4 2.93234437E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1812_885012010012_6.8nF
*******
.subckt 1812_885012010013_10nF 1 2
Rser 1 3 0.0378661246646
Lser 2 4 3.63058436E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012010013_10nF
*******
.subckt 1812_885012010014_15nF 1 2
Rser 1 3 0.0258373805332
Lser 2 4 2.604228E-10
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1812_885012010014_15nF
*******
.subckt 1812_885012010015_22nF 1 2
Rser 1 3 0.0234
Lser 2 4 0.000000001
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1812_885012010015_22nF
*******
.subckt 1812_885012010016_33nF 1 2
Rser 1 3 0.0536968994705
Lser 2 4 3.37435968E-10
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1812_885012010016_33nF
*******
.subckt 1812_885012210013_1nF 1 2
Rser 1 3 0.22122
Lser 2 4 0.00000000021688
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1812_885012210013_1nF
*******
.subckt 1812_885012210014_1.5nF 1 2
Rser 1 3 0.17474
Lser 2 4 0.00000000020664
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1812_885012210014_1.5nF
*******
.subckt 1812_885012210015_2.2nF 1 2
Rser 1 3 0.13333
Lser 2 4 0.00000000015464
C1 3 4 0.0000000022
Rpar 3 4 10000000000
.ends 1812_885012210015_2.2nF
*******
.subckt 1812_885012210016_3.3nF 1 2
Rser 1 3 0.11987
Lser 2 4 0.00000000054219
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1812_885012210016_3.3nF
*******
.subckt 1812_885012210017_4.7nF 1 2
Rser 1 3 0.08329
Lser 2 4 0.00000000014772
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1812_885012210017_4.7nF
*******
.subckt 1812_885012210018_6.8nF 1 2
Rser 1 3 0.08602
Lser 2 4 0.00000000061736
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1812_885012210018_6.8nF
*******
.subckt 1812_885012210019_10nF 1 2
Rser 1 3 0.07293
Lser 2 4 0.00000000052871
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1812_885012210019_10nF
*******
.subckt 1812_885012210020_15nF 1 2
Rser 1 3 0.067
Lser 2 4 0.0000000007302
C1 3 4 0.000000015
Rpar 3 4 10000000000
.ends 1812_885012210020_15nF
*******
.subckt 1812_885012210021_22nF 1 2
Rser 1 3 0.05662
Lser 2 4 0.00000000062074
C1 3 4 0.000000022
Rpar 3 4 10000000000
.ends 1812_885012210021_22nF
*******
.subckt 1812_885012210022_33nF 1 2
Rser 1 3 0.03888
Lser 2 4 0.00000000053993
C1 3 4 0.000000033
Rpar 3 4 10000000000
.ends 1812_885012210022_33nF
*******
.subckt 1812_885012210023_47nF 1 2
Rser 1 3 0.0333
Lser 2 4 0.00000000024107
C1 3 4 0.000000047
Rpar 3 4 10000000000
.ends 1812_885012210023_47nF
*******
.subckt 1812_885012210024_68nF 1 2
Rser 1 3 0.0283
Lser 2 4 0.00000000079079
C1 3 4 0.000000068
Rpar 3 4 7400000000
.ends 1812_885012210024_68nF
*******
.subckt 1812_885012210025_100nF 1 2
Rser 1 3 0.0434286733285
Lser 2 4 5.51116314E-10
C1 3 4 0.0000001
Rpar 3 4 5000000000
.ends 1812_885012210025_100nF
*******
.subckt 1812_885012210026_150nF 1 2
Rser 1 3 0.0274984909595
Lser 2 4 6.78013757E-10
C1 3 4 0.00000015
Rpar 3 4 3300000000
.ends 1812_885012210026_150nF
*******
.subckt 1812_885012210027_220nF 1 2
Rser 1 3 0.0210915166325
Lser 2 4 5.00831292E-10
C1 3 4 0.00000022
Rpar 3 4 2300000000
.ends 1812_885012210027_220nF
*******
.subckt 1812_885012210028_330nF 1 2
Rser 1 3 0.0146375735099
Lser 2 4 4.50409847E-10
C1 3 4 0.00000033
Rpar 3 4 1500000000
.ends 1812_885012210028_330nF
*******
.subckt 1812_885012210029_470nF 1 2
Rser 1 3 0.0117735855692
Lser 2 4 3.80795098E-10
C1 3 4 0.00000047
Rpar 3 4 1100000000
.ends 1812_885012210029_470nF
*******
.subckt 1812_885012210030_680nF 1 2
Rser 1 3 0.00705429391862
Lser 2 4 4.5048548E-10
C1 3 4 0.00000068
Rpar 3 4 700000000
.ends 1812_885012210030_680nF
*******
.subckt 1812_885012210031_1uF 1 2
Rser 1 3 0.00507618175382
Lser 2 4 5.00373592E-10
C1 3 4 0.000001
Rpar 3 4 500000000
.ends 1812_885012210031_1uF
*******
.subckt 1812_885012210032_2.2uF 1 2
Rser 1 3 0.00377371050938
Lser 2 4 4.19292053E-10
C1 3 4 0.0000022
Rpar 3 4 200000000
.ends 1812_885012210032_2.2uF
*******
.subckt 2220_885012214005_10uF 1 2
Rser 1 3 0.003
Lser 2 4 0.0000000012
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 2220_885012214005_10uF
*******
