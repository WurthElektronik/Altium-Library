**************************************************
* Manufacturer:           W�rth Elektronik
* Kinds:                  MLCCs - Multilayer Ceramic Chip Capacitors
* Matchcode:              WCAP-CSGP_6-3V
* Library Type:           LTspice
* Version:                rev25a
* Created/modified by:    Ella
* Date and Time:          5/19/2025
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2025 W�rth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While W�rth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, W�rth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does W�rth Elektronik eiSos guarantee that the simulation model is current.
* W�rth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* W�rth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 0402_885012005074_10pF 1 2
Rser 1 3 0.421651463477
Lser 2 4 4.14790783E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0402_885012005074_10pF
*******
.subckt 0402_885012005077_33pF 1 2
Rser 1 3 0.221604982314
Lser 2 4 3.49022204E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0402_885012005077_33pF
*******
.subckt 0402_885012005078_47pF 1 2
Rser 1 3 0.24210526915
Lser 2 4 4.45579658E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0402_885012005078_47pF
*******
.subckt 0402_885012005079_68pF 1 2
Rser 1 3 0.204212177962
Lser 2 4 3.70169713E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0402_885012005079_68pF
*******
.subckt 0402_885012005080_100pF 1 2
Rser 1 3 0.117553952575
Lser 2 4 3.96667338E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0402_885012005080_100pF
*******
.subckt 0402_885012005083_2.2pF 1 2
Rser 1 3 0.644
Lser 2 4 0.00000000032
C1 3 4 0.0000000000022
Rpar 3 4 10000000000
.ends 0402_885012005083_2.2pF
*******
.subckt 0402_885012005085_8.2pF 1 2
Rser 1 3 0.352598551895
Lser 2 4 4.16869039E-10
C1 3 4 0.0000000000082
Rpar 3 4 10000000000
.ends 0402_885012005085_8.2pF
*******
.subckt 0402_885012205080_1nF 1 2
Rser 1 3 0.266
Lser 2 4 0.0000000008
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0402_885012205080_1nF
*******
.subckt 0402_885012205084_4.7nF 1 2
Rser 1 3 0.155
Lser 2 4 0.0000000004
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0402_885012205084_4.7nF
*******
.subckt 0603_885012006073_10pF 1 2
Rser 1 3 0.407424144741
Lser 2 4 5.41304078E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0603_885012006073_10pF
*******
.subckt 0603_885012006074_15pF 1 2
Rser 1 3 0.380584852252
Lser 2 4 5.65804545E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0603_885012006074_15pF
*******
.subckt 0603_885012006076_33pF 1 2
Rser 1 3 0.286862998414
Lser 2 4 6.50561095E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0603_885012006076_33pF
*******
.subckt 0603_885012006077_47pF 1 2
Rser 1 3 0.245803082005
Lser 2 4 6.35972597E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0603_885012006077_47pF
*******
.subckt 0603_885012006078_68pF 1 2
Rser 1 3 0.200732636434
Lser 2 4 5.98671906E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0603_885012006078_68pF
*******
.subckt 0603_885012006079_100pF 1 2
Rser 1 3 0.147736548124
Lser 2 4 5.50713639E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012006079_100pF
*******
.subckt 0603_885012006080_150pF 1 2
Rser 1 3 0.123096464746
Lser 2 4 5.27226081E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012006080_150pF
*******
.subckt 0603_885012006082_330pF 1 2
Rser 1 3 0.0953300210797
Lser 2 4 4.24072373E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012006082_330pF
*******
.subckt 0603_885012006083_470pF 1 2
Rser 1 3 0.0701382798145
Lser 2 4 4.13398494E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012006083_470pF
*******
.subckt 0603_885012006084_680pF 1 2
Rser 1 3 0.0621072894488
Lser 2 4 4.13475086E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012006084_680pF
*******
.subckt 0603_885012006085_1nF 1 2
Rser 1 3 0.0532527583524
Lser 2 4 3.27557981E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012006085_1nF
*******
.subckt 0603_885012206102_100pF 1 2
Rser 1 3 0.903793201449
Lser 2 4 4.30927368E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0603_885012206102_100pF
*******
.subckt 0603_885012206103_150pF 1 2
Rser 1 3 0.663307587764
Lser 2 4 4.01639305E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0603_885012206103_150pF
*******
.subckt 0603_885012206105_330pF 1 2
Rser 1 3 0.471881844186
Lser 2 4 4.17174312E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0603_885012206105_330pF
*******
.subckt 0603_885012206106_470pF 1 2
Rser 1 3 0.3
Lser 2 4 0.000000000401
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0603_885012206106_470pF
*******
.subckt 0603_885012206107_680pF 1 2
Rser 1 3 0.307694453707
Lser 2 4 4.68126223E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0603_885012206107_680pF
*******
.subckt 0603_885012206108_1nF 1 2
Rser 1 3 0.202024514637
Lser 2 4 5.1469819E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0603_885012206108_1nF
*******
.subckt 0603_885012206109_1.5nF 1 2
Rser 1 3 0.160907873586
Lser 2 4 4.36594994E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0603_885012206109_1.5nF
*******
.subckt 0603_885012206111_3.3nF 1 2
Rser 1 3 0.141390340152
Lser 2 4 5.69446762E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0603_885012206111_3.3nF
*******
.subckt 0603_885012206112_4.7nF 1 2
Rser 1 3 0.0887774662878
Lser 2 4 4.3949757E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0603_885012206112_4.7nF
*******
.subckt 0603_885012206113_6.8nF 1 2
Rser 1 3 0.0566471875739
Lser 2 4 4.04270889E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0603_885012206113_6.8nF
*******
.subckt 0603_885012206114_10nF 1 2
Rser 1 3 0.0614305159536
Lser 2 4 4.58570264E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206114_10nF
*******
.subckt 0603_885012206118_47nF 1 2
Rser 1 3 0.0260966431276
Lser 2 4 4.02961106E-10
C1 3 4 0.000000047
Rpar 3 4 2100000000
.ends 0603_885012206118_47nF
*******
.subckt 0603_885012206120_100nF 1 2
Rser 1 3 0.02
Lser 2 4 0.0000000008
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0603_885012206120_100nF
*******
.subckt 0603_885012206114R_10nF 1 2
Rser 1 3 0.0614305159536
Lser 2 4 4.58570264E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0603_885012206114R_10nF
*******
.subckt 0805_885012007076_10pF 1 2
Rser 1 3 0.348978588999
Lser 2 4 4.65201661E-10
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 0805_885012007076_10pF
*******
.subckt 0805_885012007077_15pF 1 2
Rser 1 3 0.299948487506
Lser 2 4 4.54423504E-10
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 0805_885012007077_15pF
*******
.subckt 0805_885012007079_33pF 1 2
Rser 1 3 0.121980282644
Lser 2 4 4.43859848E-10
C1 3 4 0.000000000033
Rpar 3 4 10000000000
.ends 0805_885012007079_33pF
*******
.subckt 0805_885012007080_47pF 1 2
Rser 1 3 0.166811229395
Lser 2 4 4.10637959E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 0805_885012007080_47pF
*******
.subckt 0805_885012007081_68pF 1 2
Rser 1 3 0.180760159531
Lser 2 4 3.86267029E-10
C1 3 4 0.000000000068
Rpar 3 4 10000000000
.ends 0805_885012007081_68pF
*******
.subckt 0805_885012007082_100pF 1 2
Rser 1 3 0.0753079048439
Lser 2 4 2.90973988E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012007082_100pF
*******
.subckt 0805_885012007083_150pF 1 2
Rser 1 3 0.198942265358
Lser 2 4 3.89898948E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012007083_150pF
*******
.subckt 0805_885012007085_330pF 1 2
Rser 1 3 0.0776936134254
Lser 2 4 2.60803415E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012007085_330pF
*******
.subckt 0805_885012007086_470pF 1 2
Rser 1 3 0.0588553647502
Lser 2 4 2.97840521E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012007086_470pF
*******
.subckt 0805_885012007087_680pF 1 2
Rser 1 3 0.0627822674091
Lser 2 4 2.56856486E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012007087_680pF
*******
.subckt 0805_885012007088_1nF 1 2
Rser 1 3 0.0369190815603
Lser 2 4 3.02824205E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012007088_1nF
*******
.subckt 0805_885012007089_1.5nF 1 2
Rser 1 3 0.0444913409463
Lser 2 4 3.70041338E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012007089_1.5nF
*******
.subckt 0805_885012007091_3.3nF 1 2
Rser 1 3 0.0238862333296
Lser 2 4 3.52340361E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012007091_3.3nF
*******
.subckt 0805_885012007092_4.7nF 1 2
Rser 1 3 0.0360290329923
Lser 2 4 3.13853583E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012007092_4.7nF
*******
.subckt 0805_885012207110_100pF 1 2
Rser 1 3 0.893542107954
Lser 2 4 3.72840309E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 0805_885012207110_100pF
*******
.subckt 0805_885012207111_150pF 1 2
Rser 1 3 0.75393192763
Lser 2 4 4.30786527E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 0805_885012207111_150pF
*******
.subckt 0805_885012207113_330pF 1 2
Rser 1 3 0.884149804092
Lser 2 4 3.16830341E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 0805_885012207113_330pF
*******
.subckt 0805_885012207114_470pF 1 2
Rser 1 3 0.374236748173
Lser 2 4 4.69987959E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 0805_885012207114_470pF
*******
.subckt 0805_885012207115_680pF 1 2
Rser 1 3 0.441399652418
Lser 2 4 3.85533833E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 0805_885012207115_680pF
*******
.subckt 0805_885012207116_1nF 1 2
Rser 1 3 0.200201288389
Lser 2 4 4.27706413E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 0805_885012207116_1nF
*******
.subckt 0805_885012207117_1.5nF 1 2
Rser 1 3 0.165813253283
Lser 2 4 4.70069305E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 0805_885012207117_1.5nF
*******
.subckt 0805_885012207119_3.3nF 1 2
Rser 1 3 0.107994017051
Lser 2 4 4.67027278E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 0805_885012207119_3.3nF
*******
.subckt 0805_885012207120_4.7nF 1 2
Rser 1 3 0.0819387083384
Lser 2 4 4.01268553E-10
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 0805_885012207120_4.7nF
*******
.subckt 0805_885012207121_6.8nF 1 2
Rser 1 3 0.0730376666068
Lser 2 4 4.71078792E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 0805_885012207121_6.8nF
*******
.subckt 0805_885012207122_10nF 1 2
Rser 1 3 0.0602542793423
Lser 2 4 5.20580851E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 0805_885012207122_10nF
*******
.subckt 0805_885012207123_15nF 1 2
Rser 1 3 0.0418698831686
Lser 2 4 4.51086218E-10
C1 3 4 0.000000015
Rpar 3 4 6700000000
.ends 0805_885012207123_15nF
*******
.subckt 0805_885012207124_22nF 1 2
Rser 1 3 0.05
Lser 2 4 5.34340678E-10
C1 3 4 0.000000022
Rpar 3 4 4500000000
.ends 0805_885012207124_22nF
*******
.subckt 0805_885012207125_33nF 1 2
Rser 1 3 0.027855481442
Lser 2 4 4.0266816E-10
C1 3 4 0.000000033
Rpar 3 4 3000000000
.ends 0805_885012207125_33nF
*******
.subckt 0805_885012207126_47nF 1 2
Rser 1 3 0.0193681345947
Lser 2 4 3.56511593E-10
C1 3 4 0.000000047
Rpar 3 4 2100000000
.ends 0805_885012207126_47nF
*******
.subckt 0805_885012207127_68nF 1 2
Rser 1 3 0.0131992658565
Lser 2 4 3.66797021E-10
C1 3 4 0.000000068
Rpar 3 4 1500000000
.ends 0805_885012207127_68nF
*******
.subckt 0805_885012207128_100nF 1 2
Rser 1 3 0.0114794409661
Lser 2 4 3.71233852E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 0805_885012207128_100nF
*******
.subckt 0805_885012207130_470nF 1 2
Rser 1 3 0.011
Lser 2 4 0.0000000009
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 0805_885012207130_470nF
*******
.subckt 1206_885012008061_10pF 1 2
Rser 1 3 0.3685
Lser 2 4 0.00000000065
C1 3 4 0.00000000001
Rpar 3 4 10000000000
.ends 1206_885012008061_10pF
*******
.subckt 1206_885012008062_15pF 1 2
Rser 1 3 0.35
Lser 2 4 0.00000000056
C1 3 4 0.000000000015
Rpar 3 4 10000000000
.ends 1206_885012008062_15pF
*******
.subckt 1206_885012008065_47pF 1 2
Rser 1 3 0.19407783985
Lser 2 4 5.43052823E-10
C1 3 4 0.000000000047
Rpar 3 4 10000000000
.ends 1206_885012008065_47pF
*******
.subckt 1206_885012008067_100pF 1 2
Rser 1 3 0.157459451422
Lser 2 4 4.64194319E-10
C1 3 4 0.0000000001
Rpar 3 4 10000000000
.ends 1206_885012008067_100pF
*******
.subckt 1206_885012008068_150pF 1 2
Rser 1 3 0.130548247324
Lser 2 4 4.36494773E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012008068_150pF
*******
.subckt 1206_885012008070_330pF 1 2
Rser 1 3 0.0931468259828
Lser 2 4 4.33607632E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012008070_330pF
*******
.subckt 1206_885012008071_470pF 1 2
Rser 1 3 0.0863181912042
Lser 2 4 4.5763957E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012008071_470pF
*******
.subckt 1206_885012008072_680pF 1 2
Rser 1 3 0.0777497909642
Lser 2 4 4.75215911E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012008072_680pF
*******
.subckt 1206_885012008073_1nF 1 2
Rser 1 3 0.0477152917275
Lser 2 4 4.99751981E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012008073_1nF
*******
.subckt 1206_885012008074_1.5nF 1 2
Rser 1 3 0.0354598757287
Lser 2 4 3.99445906E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012008074_1.5nF
*******
.subckt 1206_885012008076_3.3nF 1 2
Rser 1 3 0.0314389546323
Lser 2 4 4.34527012E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012008076_3.3nF
*******
.subckt 1206_885012008078_6.8nF 1 2
Rser 1 3 0.0257323206072
Lser 2 4 4.35781903E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012008078_6.8nF
*******
.subckt 1206_885012008079_10nF 1 2
Rser 1 3 0.0235458917441
Lser 2 4 4.56933086E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012008079_10nF
*******
.subckt 1206_885012208101_150pF 1 2
Rser 1 3 0.70365102611
Lser 2 4 3.78992769E-10
C1 3 4 0.00000000015
Rpar 3 4 10000000000
.ends 1206_885012208101_150pF
*******
.subckt 1206_885012208103_330pF 1 2
Rser 1 3 0.416289638796
Lser 2 4 4.89828253E-10
C1 3 4 0.00000000033
Rpar 3 4 10000000000
.ends 1206_885012208103_330pF
*******
.subckt 1206_885012208104_470pF 1 2
Rser 1 3 0.362109688542
Lser 2 4 4.01551911E-10
C1 3 4 0.00000000047
Rpar 3 4 10000000000
.ends 1206_885012208104_470pF
*******
.subckt 1206_885012208105_680pF 1 2
Rser 1 3 0.332767276854
Lser 2 4 5.5598151E-10
C1 3 4 0.00000000068
Rpar 3 4 10000000000
.ends 1206_885012208105_680pF
*******
.subckt 1206_885012208106_1nF 1 2
Rser 1 3 0.24361864545
Lser 2 4 4.48764151E-10
C1 3 4 0.000000001
Rpar 3 4 10000000000
.ends 1206_885012208106_1nF
*******
.subckt 1206_885012208107_1.5nF 1 2
Rser 1 3 0.185507432166
Lser 2 4 4.5702585E-10
C1 3 4 0.0000000015
Rpar 3 4 10000000000
.ends 1206_885012208107_1.5nF
*******
.subckt 1206_885012208109_3.3nF 1 2
Rser 1 3 0.123971561911
Lser 2 4 4.87780525E-10
C1 3 4 0.0000000033
Rpar 3 4 10000000000
.ends 1206_885012208109_3.3nF
*******
.subckt 1206_885012208110_4.7nF 1 2
Rser 1 3 0.1
Lser 2 4 0.00000000049
C1 3 4 0.0000000047
Rpar 3 4 10000000000
.ends 1206_885012208110_4.7nF
*******
.subckt 1206_885012208111_6.8nF 1 2
Rser 1 3 0.0785959830702
Lser 2 4 5.43016322E-10
C1 3 4 0.0000000068
Rpar 3 4 10000000000
.ends 1206_885012208111_6.8nF
*******
.subckt 1206_885012208112_10nF 1 2
Rser 1 3 0.0821267479008
Lser 2 4 5.05894889E-10
C1 3 4 0.00000001
Rpar 3 4 10000000000
.ends 1206_885012208112_10nF
*******
.subckt 1206_885012208113_15nF 1 2
Rser 1 3 0.0562607370369
Lser 2 4 5.19798206E-10
C1 3 4 0.000000015
Rpar 3 4 6700000000
.ends 1206_885012208113_15nF
*******
.subckt 1206_885012208115_33nF 1 2
Rser 1 3 0.0633889215043
Lser 2 4 5.17142938E-10
C1 3 4 0.000000033
Rpar 3 4 3000000000
.ends 1206_885012208115_33nF
*******
.subckt 1206_885012208116_47nF 1 2
Rser 1 3 0.0362676531527
Lser 2 4 5.26289035E-10
C1 3 4 0.000000047
Rpar 3 4 2100000000
.ends 1206_885012208116_47nF
*******
.subckt 1206_885012208117_68nF 1 2
Rser 1 3 0.0206252921491
Lser 2 4 4.8689903E-10
C1 3 4 0.000000068
Rpar 3 4 1500000000
.ends 1206_885012208117_68nF
*******
.subckt 1206_885012208118_100nF 1 2
Rser 1 3 0.0147498855833
Lser 2 4 5.50636098E-10
C1 3 4 0.0000001
Rpar 3 4 1000000000
.ends 1206_885012208118_100nF
*******
.subckt 1206_885012208119_150nF 1 2
Rser 1 3 0.00800974723287
Lser 2 4 3.65669763E-10
C1 3 4 0.00000015
Rpar 3 4 700000000
.ends 1206_885012208119_150nF
*******
.subckt 1206_885012208122_470nF 1 2
Rser 1 3 0.010704092868
Lser 2 4 6.6200966E-10
C1 3 4 0.00000047
Rpar 3 4 200000000
.ends 1206_885012208122_470nF
*******
.subckt 1206_885012208124_2.2uF 1 2
Rser 1 3 0.015
Lser 2 4 0.0000000030781
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 1206_885012208124_2.2uF
*******
.subckt 1210_885012209069_1uF 1 2
Rser 1 3 0.0053441098735
Lser 2 4 6.51295361E-10
C1 3 4 0.000001
Rpar 3 4 100000000
.ends 1210_885012209069_1uF
*******
.subckt 1210_885012209071_2.2uF 1 2
Rser 1 3 0.014
Lser 2 4 0.000000000755
C1 3 4 0.0000022
Rpar 3 4 50000000
.ends 1210_885012209071_2.2uF
*******
.subckt 2220_885012214002_3.3uF 1 2
Rser 1 3 0.0056
Lser 2 4 0.0000000012
C1 3 4 0.0000033
Rpar 3 4 30000000
.ends 2220_885012214002_3.3uF
*******
.subckt 2220_885012214003_4.7uF 1 2
Rser 1 3 0.0043
Lser 2 4 0.0000000013
C1 3 4 0.0000047
Rpar 3 4 20000000
.ends 2220_885012214003_4.7uF
*******
.subckt 2220_885012214001_10uF 1 2
Rser 1 3 0.003
Lser 2 4 0.0000000012
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 2220_885012214001_10uF
*******
.subckt 2220_885012214006_10uF 1 2
Rser 1 3 0.003
Lser 2 4 0.0000000012
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 2220_885012214006_10uF
*******
