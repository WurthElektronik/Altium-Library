**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  High Frequency SMT Inductor
* Matchcode:              WE-GFH 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-09
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 2520_7447629010_1u 1 2
Rp 1 2 4462
Cp 1 2 0.277p
Rs 1 N3 0.34
L1 N3 2 0.957u
.ends 2520_7447629010_1u
*******
.subckt 2520_7447629015_1.5u 1 2
Rp 1 2 2845.86
Cp 1 2 0.961p
Rs 1 N3 0.393
L1 N3 2 1.5u
.ends 2520_7447629015_1.5u
*******
.subckt 2520_7447629022_2.2u 1 2
Rp 1 2 3345.25
Cp 1 2 1.827p
Rs 1 N3 0.51
L1 N3 2 2.2u
.ends 2520_7447629022_2.2u
*******
.subckt 2520_7447629033_3.3u 1 2
Rp 1 2 4676.71
Cp 1 2 2.251p
Rs 1 N3 0.625
L1 N3 2 3.3u
.ends 2520_7447629033_3.3u
*******
.subckt 2520_7447629047_4.7u 1 2
Rp 1 2 5593.74
Cp 1 2 2.203p
Rs 1 N3 0.75
L1 N3 2 4.7u
.ends 2520_7447629047_4.7u
*******
.subckt 2520_7447629068_6.8u 1 2
Rp 1 2 7706.21
Cp 1 2 2.091p
Rs 1 N3 0.96
L1 N3 2 6.8u
.ends 2520_7447629068_6.8u
*******
.subckt 2520_7447629100_10u 1 2
Rp 1 2 9172.38
Cp 1 2 2.842p
Rs 1 N3 1.7
L1 N3 2 10u
.ends 2520_7447629100_10u
*******
.subckt 2520_7447629150_15u 1 2
Rp 1 2 12435.4
Cp 1 2 3.285p
Rs 1 N3 2.11
L1 N3 2 15u
.ends 2520_7447629150_15u
*******
.subckt 2520_7447629220_22u 1 2
Rp 1 2 16159.7
Cp 1 2 2.85p
Rs 1 N3 2.762
L1 N3 2 22u
.ends 2520_7447629220_22u
*******
.subckt 2520_7447629330_33u 1 2
Rp 1 2 21163
Cp 1 2 3.208p
Rs 1 N3 4.3
L1 N3 2 33u
.ends 2520_7447629330_33u
*******
.subckt 3225_744764901_1u 1 2
Rp 1 2 2887.58
Cp 1 2 0.706p
Rs 1 N3 0.14
L1 N3 2 1u
.ends 3225_744764901_1u
*******
.subckt 3225_7447649015_1.5u 1 2
Rp 1 2 3790
Cp 1 2 1.24p
Rs 1 N3 0.17
L1 N3 2 1.49u
.ends 3225_7447649015_1.5u
*******
.subckt 3225_744764902_2.2u 1 2
Rp 1 2 6355.45
Cp 1 2 1.24p
Rs 1 N3 0.234
L1 N3 2 2.2u
.ends 3225_744764902_2.2u
*******
.subckt 3225_744764903_3.3u 1 2
Rp 1 2 7525.99
Cp 1 2 1.357p
Rs 1 N3 0.293
L1 N3 2 3.3u
.ends 3225_744764903_3.3u
*******
.subckt 3225_744764904_4.7u 1 2
Rp 1 2 9543.57
Cp 1 2 1.389p
Rs 1 N3 0.468
L1 N3 2 4.7u
.ends 3225_744764904_4.7u
*******
.subckt 3225_744764910_10u 1 2
Rp 1 2 15035
Cp 1 2 1397p
Rs 1 N3 1
L1 N3 2 9.9u
.ends 3225_744764910_10u
*******
.subckt 3225_7447649115_15u 1 2
Rp 1 2 20192
Cp 1 2 1.298p
Rs 1 N3 1.521
L1 N3 2 15.57u
.ends 3225_7447649115_15u
*******
.subckt 3225_7447649122_22u 1 2
Rp 1 2 28531.3
Cp 1 2 1.553p
Rs 1 N3 2.34
L1 N3 2 22u
.ends 3225_7447649122_22u
*******
.subckt 3225_7447649133_33u 1 2
Rp 1 2 38263.3
Cp 1 2 1.707p
Rs 1 N3 3.276
L1 N3 2 33u
.ends 3225_7447649133_33u
*******
.subckt 3225_7447649147_47u 1 2
Rp 1 2 43978
Cp 1 2 1.49p
Rs 1 N3 4.914
L1 N3 2 46.027u
.ends 3225_7447649147_47u
*******
.subckt 3225_7447649168_68u 1 2
Rp 1 2 188392
Cp 1 2 1.789p
Rs 1 N3 7.605
L1 N3 2 68u
.ends 3225_7447649168_68u
*******
.subckt 3225_744764920_100u 1 2
Rp 1 2 76383.9
Cp 1 2 1.692p
Rs 1 N3 9.126
L1 N3 2 100u
.ends 3225_744764920_100u
*******
.subckt 4532_744766901_1u 1 2
Rp 1 2 3105.29
Cp 1 2 0.438p
Rs 1 N3 0.081
L1 N3 2 1u
.ends 4532_744766901_1u
*******
.subckt 4532_7447669012_1.2u 1 2
Rp 1 2 3727.35
Cp 1 2 0.747p
Rs 1 N3 0.093
L1 N3 2 1.2u
.ends 4532_7447669012_1.2u
*******
.subckt 4532_744766902_2.2u 1 2
Rp 1 2 4089
Cp 1 2 1.738p
Rs 1 N3 0.144
L1 N3 2 2.159u
.ends 4532_744766902_2.2u
*******
.subckt 4532_744766903_3.3u 1 2
Rp 1 2 6617.99
Cp 1 2 2.342p
Rs 1 N3 0.178
L1 N3 2 3.3u
.ends 4532_744766903_3.3u
*******
.subckt 4532_7447669039_3.9u 1 2
Rp 1 2 7957
Cp 1 2 1.93p
Rs 1 N3 0.2
L1 N3 2 3.785u
.ends 4532_7447669039_3.9u
*******
.subckt 4532_744766904_4.7u 1 2
Rp 1 2 7628.48
Cp 1 2 2.096p
Rs 1 N3 0.215
L1 N3 2 4.7u
.ends 4532_744766904_4.7u
*******
.subckt 4532_744766906_6.8u 1 2
Rp 1 2 13363.8
Cp 1 2 2.32p
Rs 1 N3 0.271
L1 N3 2 6.8u
.ends 4532_744766906_6.8u
*******
.subckt 4532_744766910_10u 1 2
Rp 1 2 18622
Cp 1 2 2.091p
Rs 1 N3 0.405
L1 N3 2 10u
.ends 4532_744766910_10u
*******
.subckt 4532_7447669112_12u 1 2
Rp 1 2 20890.6
Cp 1 2 2.343p
Rs 1 N3 0.444
L1 N3 2 12u
.ends 4532_7447669112_12u
*******
.subckt 4532_7447669115_15u 1 2
Rp 1 2 24670.2
Cp 1 2 2.499p
Rs 1 N3 0.511
L1 N3 2 15u
.ends 4532_7447669115_15u
*******
.subckt 4532_7447669118_18u 1 2
Rp 1 2 32480.2
Cp 1 2 2.479p
Rs 1 N3 0.654
L1 N3 2 18u
.ends 4532_7447669118_18u
*******
.subckt 4532_7447669122_22u 1 2
Rp 1 2 42816.1
Cp 1 2 2.252p
Rs 1 N3 0.767
L1 N3 2 22u
.ends 4532_7447669122_22u
*******
.subckt 4532_7447669127_27u 1 2
Rp 1 2 44704.7
Cp 1 2 2.494p
Rs 1 N3 0.849
L1 N3 2 27u
.ends 4532_7447669127_27u
*******
.subckt 4532_7447669133_33u 1 2
Rp 1 2 38959
Cp 1 2 2.331p
Rs 1 N3 1.4
L1 N3 2 33.045u
.ends 4532_7447669133_33u
*******
.subckt 4532_7447669139_39u 1 2
Rp 1 2 35992
Cp 1 2 2.127p
Rs 1 N3 1.6
L1 N3 2 38.785u
.ends 4532_7447669139_39u
*******
.subckt 4532_7447669147_47u 1 2
Rp 1 2 91375.1
Cp 1 2 2.349p
Rs 1 N3 1.46
L1 N3 2 47u
.ends 4532_7447669147_47u
*******
.subckt 4532_7447669156_56u 1 2
Rp 1 2 133478
Cp 1 2 2.449p
Rs 1 N3 1.94
L1 N3 2 56u
.ends 4532_7447669156_56u
*******
.subckt 4532_7447669168_68u 1 2
Rp 1 2 144173
Cp 1 2 2.585p
Rs 1 N3 2.195
L1 N3 2 68u
.ends 4532_7447669168_68u
*******
.subckt 4532_7447669182_82u 1 2
Rp 1 2 256010
Cp 1 2 2.572p
Rs 1 N3 3.11
L1 N3 2 82u
.ends 4532_7447669182_82u
*******
.subckt 4532_744766920_100u 1 2
Rp 1 2 317330
Cp 1 2 2.454p
Rs 1 N3 3.56
L1 N3 2 100u
.ends 4532_744766920_100u
*******
.subckt 4532_7447669212_120u 1 2
Rp 1 2 476140
Cp 1 2 2.417p
Rs 1 N3 4.185
L1 N3 2 120u
.ends 4532_7447669212_120u
*******
.subckt 4532_7447669218_180u 1 2
Rp 1 2 277120
Cp 1 2 2.612p
Rs 1 N3 6.15
L1 N3 2 180u
.ends 4532_7447669218_180u
*******
.subckt 4532_7447669220_220u 1 2
Rp 1 2 188174
Cp 1 2 2.309p
Rs 1 N3 6.94
L1 N3 2 220u
.ends 4532_7447669220_220u
*******
