**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT EMI Suppression Ferrite Bead
* Matchcode:             WE-CBA
* Library Type:          LTspice
* Version:               rev21a
* Created/modified by:   Ella
* Date and Time:         2022/11/4
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
.subckt 0201_782219100_10ohm 1 2
Rp 1 2 14.001647
Cp 1 2 1.31p
Rs 1 N3 0.055
L1 N3 2 0.020856937u
.ends 0201_782219100_10ohm
*******
.subckt 0201_782219600_60ohm 1 2
Rp 1 2 127.679039
Cp 1 2 0.138786005p
Rs 1 N3 0.25
L1 N3 2 0.098234695u
.ends 0201_782219600_60ohm
*******
.subckt 0201_782219121_120ohm 1 2
Rp 1 2 157.473156
Cp 1 2 0.303648583p
Rs 1 N3 0.29
L1 N3 2 0.266321573u
.ends 0201_782219121_120ohm
*******
.subckt 0201_782219241_240ohm 1 2
Rp 1 2 377.648044
Cp 1 2 0.385147298p
Rs 1 N3 0.57
L1 N3 2 0.462853473u
.ends 0201_782219241_240ohm
*******
.subckt 0201_782219301_300ohm 1 2
Rp 1 2 499.785512
Cp 1 2 0.341711468p
Rs 1 N3 0.61
L1 N3 2 0.556682313u
.ends 0201_782219301_300ohm
*******
.subckt 0201_782219561_560ohm 1 2
Rp 1 2 788.750819
Cp 1 2 0.55p
Rs 1 N3 0.75
L1 N3 2 1.747131u
.ends 0201_782219561_560ohm
*******
.subckt 0402_782422101_100ohm 1 2
Rp 1 2 120.5
Cp 1 2 0.279p
Rs 1 N3 0.3
L1 N3 2 0.6u
.ends 0402_782422101_100ohm
*******
.subckt 0402_782422102_1000ohm 1 2
Rp 1 2 1050
Cp 1 2 0.59p
Rs 1 N3 1
L1 N3 2 1.8u
.ends 0402_782422102_1000ohm
*******
.subckt 0402_782422121_120ohm 1 2
Rp 1 2 182
Cp 1 2 0.343p
Rs 1 N3 0.2
L1 N3 2 0.505u
.ends 0402_782422121_120ohm
*******
.subckt 0402_782422181_180ohm 1 2
Rp 1 2 230
Cp 1 2 0.288p
Rs 1 N3 0.3
L1 N3 2 0.39u
.ends 0402_782422181_180ohm
*******
.subckt 0402_782422221_220ohm 1 2
Rp 1 2 330
Cp 1 2 0.37p
Rs 1 N3 0.3
L1 N3 2 0.43u
.ends 0402_782422221_220ohm
*******
.subckt 0402_782422231_220ohm 1 2
Rp 1 2 270
Cp 1 2 0.42p
Rs 1 N3 0.35
L1 N3 2 0.67u
.ends 0402_782422231_220ohm
*******
.subckt 0402_782422241_240ohm 1 2
Rp 1 2 361
Cp 1 2 0.275p
Rs 1 N3 0.35
L1 N3 2 0.911u
.ends 0402_782422241_240ohm
*******
.subckt 0402_782422301_300ohm 1 2
Rp 1 2 332
Cp 1 2 0.316p
Rs 1 N3 0.7
L1 N3 2 0.076u
.ends 0402_782422301_300ohm
*******
.subckt 0402_782422331_330ohm 1 2
Rp 1 2 535
Cp 1 2 0.445p
Rs 1 N3 0.5
L1 N3 2 0.78u
.ends 0402_782422331_330ohm
*******
.subckt 0402_782422511_510ohm 1 2
Rp 1 2 650
Cp 1 2 0.33p
Rs 1 N3 0.8
L1 N3 2 1.7u
.ends 0402_782422511_510ohm
*******
.subckt 0402_782422601_600ohm 1 2
Rp 1 2 750
Cp 1 2 0.35p
Rs 1 N3 0.8
L1 N3 2 1u
.ends 0402_782422601_600ohm
*******
.subckt 0402_782422611_600ohm 1 2
Rp 1 2 570
Cp 1 2 0.36p
Rs 1 N3 0.6
L1 N3 2 1.6u
.ends 0402_782422611_600ohm
*******
.subckt 0402_782423100_10ohm 1 2
Rp 1 2 14
Cp 1 2 0.057p
Rs 1 N3 0.03
L1 N3 2 0.0232u
.ends 0402_782423100_10ohm
*******
.subckt 0402_782423700_70ohm 1 2
Rp 1 2 154
Cp 1 2 0.349p
Rs 1 N3 0.09
L1 N3 2 0.125u
.ends 0402_782423700_70ohm
*******
.subckt 0402_782429102_1000ohm 1 2
Rp 1 2 1205.835
Cp 1 2 0.673096327p
Rs 1 N3 0.43
L1 N3 2 2.445964u
.ends 0402_782429102_1000ohm
*******
.subckt 0402_782429152_1500ohm 1 2
Rp 1 2 1533
Cp 1 2 0.623995609p
Rs 1 N3 0.43
L1 N3 2 3u
.ends 0402_782429152_1500ohm
*******
.subckt 0402_782429601_600ohm 1 2
Rp 1 2 730.563277
Cp 1 2 0.648453724p
Rs 1 N3 0.22
L1 N3 2 1.01986u
.ends 0402_782429601_600ohm
*******
.subckt 0402_782429111_110ohm 1 2
Rp 1 2 201.584103
Cp 1 2 0.4p
Rs 1 N3 0.07
L1 N3 2 0.213456094u
.ends 0402_782429111_110ohm
*******
.subckt 0402_782429161_160ohm 1 2
Rp 1 2 308.89489
Cp 1 2 0.46003571p
Rs 1 N3 0.12
L1 N3 2 0.433467564u
.ends 0402_782429161_160ohm
*******
.subckt 0402_782429261_260ohm 1 2
Rp 1 2 393.732923
Cp 1 2 0.6121285421p
Rs 1 N3 0.12
L1 N3 2 0.617816383u
.ends 0402_782429261_260ohm
*******
.subckt 0402_782429461_460ohm 1 2
Rp 1 2 1260.241
Cp 1 2 0.687046214p
Rs 1 N3 0.35
L1 N3 2 0.728916363u
.ends 0402_782429461_460ohm
*******
.subckt 0402_782429182_1800ohm 1 2
Rp 1 2 2726.742
Cp 1 2 0.053399989p
Rs 1 N3 1.91
L1 N3 2 3.050897u
.ends 0402_782429182_1800ohm
*******
.subckt 0603_782631101_100ohm 1 2
Rp 1 2 612
Cp 1 2 0.65p
Rs 1 N3 0.2
L1 N3 2 0.215u
.ends 0603_782631101_100ohm
*******
.subckt 0603_782631111_100ohm 1 2
Rp 1 2 120
Cp 1 2 0.68p
Rs 1 N3 0.12
L1 N3 2 0.034u
.ends 0603_782631111_100ohm
*******
.subckt 0603_782631131_120ohm 1 2
Rp 1 2 172
Cp 1 2 0.545p
Rs 1 N3 0.12
L1 N3 2 0.37u
.ends 0603_782631131_120ohm
*******
.subckt 0603_782631141_120ohm 1 2
Rp 1 2 140
Cp 1 2 0.56p
Rs 1 N3 0.05
L1 N3 2 0.325u
.ends 0603_782631141_120ohm
*******
.subckt 0603_782631182_1800ohm 1 2
Rp 1 2 2250
Cp 1 2 0.8p
Rs 1 N3 0.75
L1 N3 2 1.9u
.ends 0603_782631182_1800ohm
*******
.subckt 0603_782631222_2200ohm 1 2
Rp 1 2 2286
Cp 1 2 1.057p
Rs 1 N3 0.8
L1 N3 2 1.5u
.ends 0603_782631222_2200ohm
*******
.subckt 0603_782631331_330ohm 1 2
Rp 1 2 690
Cp 1 2 0.62p
Rs 1 N3 0.25
L1 N3 2 0.57u
.ends 0603_782631331_330ohm
*******
.subckt 0603_782632102_1000ohm 1 2
Rp 1 2 850
Cp 1 2 0.88p
Rs 1 N3 0.5
L1 N3 2 3.5u
.ends 0603_782632102_1000ohm
*******
.subckt 0603_782632121_120ohm 1 2
Rp 1 2 180
Cp 1 2 0.45p
Rs 1 N3 0.2
L1 N3 2 0.45u
.ends 0603_782632121_120ohm
*******
.subckt 0603_782632181_180ohm 1 2
Rp 1 2 255
Cp 1 2 0.53p
Rs 1 N3 0.2
L1 N3 2 0.5u
.ends 0603_782632181_180ohm
*******
.subckt 0603_782632511_510ohm 1 2
Rp 1 2 638
Cp 1 2 0.6p
Rs 1 N3 0.35
L1 N3 2 1.4u
.ends 0603_782632511_510ohm
*******
.subckt 0603_782632620_62ohm 1 2
Rp 1 2 90
Cp 1 2 0.64p
Rs 1 N3 0.15
L1 N3 2 0.14u
.ends 0603_782632620_62ohm
*******
.subckt 0603_782633601_600ohm 1 2
Rp 1 2 605
Cp 1 2 1.1p
Rs 1 N3 0.2
L1 N3 2 2.5u
.ends 0603_782633601_600ohm
*******
.subckt 0603_782633620_62ohm 1 2
Rp 1 2 90
Cp 1 2 0.6p
Rs 1 N3 0.04
L1 N3 2 0.21u
.ends 0603_782633620_62ohm
*******
.subckt 0603_782639220_22ohm 1 2
Rp 1 2 40
Cp 1 2 0.243p
Rs 1 N3 0.00295
L1 N3 2 0.035u
.ends 0603_782639220_22ohm
*******
.subckt 0603_782639601_600ohm 1 2
Rp 1 2 635.759722
Cp 1 2 0.83595329p
Rs 1 N3 0.09
L1 N3 2 1.000069u
.ends 0603_782639601_600ohm
*******
.subckt 0805_782851102_1000ohm 1 2
Rp 1 2 1035
Cp 1 2 1.005p
Rs 1 N3 0.35
L1 N3 2 1.08u
.ends 0805_782851102_1000ohm
*******
.subckt 0805_782851202_2200ohm 1 2
Rp 1 2 2350
Cp 1 2 0.915p
Rs 1 N3 0.45
L1 N3 2 2.25u
.ends 0805_782851202_2200ohm
*******
.subckt 0805_782851212_2000ohm 1 2
Rp 1 2 1800
Cp 1 2 0.886p
Rs 1 N3 0.42
L1 N3 2 2.6u
.ends 0805_782851212_2000ohm
*******
.subckt 0805_782853102_1000ohm 1 2
Rp 1 2 1080
Cp 1 2 1.3p
Rs 1 N3 0.3
L1 N3 2 5.3u
.ends 0805_782853102_1000ohm
*******
.subckt 0805_782853112_1100ohm 1 2
Rp 1 2 1400
Cp 1 2 1.1p
Rs 1 N3 0.3
L1 N3 2 5u
.ends 0805_782853112_1100ohm
*******
.subckt 0805_782853121_120ohm 1 2
Rp 1 2 198
Cp 1 2 1.1p
Rs 1 N3 0.035
L1 N3 2 0.38u
.ends 0805_782853121_120ohm
*******
.subckt 0805_782853131_120ohm 1 2
Rp 1 2 177
Cp 1 2 0.847p
Rs 1 N3 0.03
L1 N3 2 0.377u
.ends 0805_782853131_120ohm
*******
.subckt 0805_782853152_1500ohm 1 2
Rp 1 2 1650
Cp 1 2 1p
Rs 1 N3 0.35
L1 N3 2 6u
.ends 0805_782853152_1500ohm
*******
.subckt 0805_782853162_1500ohm 1 2
Rp 1 2 1570
Cp 1 2 1.34p
Rs 1 N3 0.3
L1 N3 2 8.3u
.ends 0805_782853162_1500ohm
*******
.subckt 0805_782853200_20ohm 1 2
Rp 1 2 33
Cp 1 2 1p
Rs 1 N3 0.008
L1 N3 2 0.05u
.ends 0805_782853200_20ohm
*******
.subckt 0805_782853221_220ohm 1 2
Rp 1 2 220
Cp 1 2 1.1p
Rs 1 N3 0.05
L1 N3 2 0.63u
.ends 0805_782853221_220ohm
*******
.subckt 0805_782853231_220ohm 1 2
Rp 1 2 360
Cp 1 2 0.68p
Rs 1 N3 0.05
L1 N3 2 0.564u
.ends 0805_782853231_220ohm
*******
.subckt 0805_782853270_27ohm 1 2
Rp 1 2 38
Cp 1 2 0.052p
Rs 1 N3 0.015
L1 N3 2 0.083u
.ends 0805_782853270_27ohm
*******
.subckt 0805_782853301_300ohm 1 2
Rp 1 2 330
Cp 1 2 1.12p
Rs 1 N3 0.05
L1 N3 2 1.21u
.ends 0805_782853301_300ohm
*******
.subckt 0805_782853321_320ohm 1 2
Rp 1 2 576.626
Cp 1 2 1.04955297286p
Rs 1 N3 0.05
L1 N3 2 0.00165041562294u
.ends 0805_782853321_320ohm
*******
.subckt 0805_782853331_330ohm 1 2
Rp 1 2 362
Cp 1 2 0.863p
Rs 1 N3 0.05
L1 N3 2 0.775u
.ends 0805_782853331_330ohm
*******
.subckt 0805_782853401_400ohm 1 2
Rp 1 2 495
Cp 1 2 1.25p
Rs 1 N3 0.3
L1 N3 2 2.07u
.ends 0805_782853401_400ohm
*******
.subckt 0805_782853561_560ohm 1 2
Rp 1 2 500
Cp 1 2 1p
Rs 1 N3 0.1
L1 N3 2 2.2u
.ends 0805_782853561_560ohm
*******
.subckt 0805_782853601_600ohm 1 2
Rp 1 2 754
Cp 1 2 0.784p
Rs 1 N3 0.3
L1 N3 2 1.381u
.ends 0805_782853601_600ohm
*******
.subckt 0805_782853611_600ohm 1 2
Rp 1 2 830
Cp 1 2 0.836p
Rs 1 N3 0.11
L1 N3 2 1.43u
.ends 0805_782853611_600ohm
*******
.subckt 0805_782853680_68ohm 1 2
Rp 1 2 110
Cp 1 2 0.83p
Rs 1 N3 0.025
L1 N3 2 0.23u
.ends 0805_782853680_68ohm
*******
.subckt 0805_782853701_700ohm 1 2
Rp 1 2 622.642880647433
Cp 1 2 1.061633380212p
Rs 1 N3 0.1
L1 N3 2 2.24477477199633E-03u
.ends 0805_782853701_700ohm
*******
.subckt 0805_782853910_91ohm 1 2
Rp 1 2 105
Cp 1 2 0.814p
Rs 1 N3 0.06
L1 N3 2 0.241u
.ends 0805_782853910_91ohm
*******
.subckt 1206_782762301_300ohm 1 2
Rp 1 2 360
Cp 1 2 1.3p
Rs 1 N3 0.1
L1 N3 2 0.95u
.ends 1206_782762301_300ohm
*******
.subckt 1206_782763102_1000ohm 1 2
Rp 1 2 1100
Cp 1 2 1.15p
Rs 1 N3 0.3
L1 N3 2 3.7u
.ends 1206_782763102_1000ohm
*******
.subckt 1206_782763301_300ohm 1 2
Rp 1 2 290
Cp 1 2 1.45p
Rs 1 N3 0.06
L1 N3 2 0.95u
.ends 1206_782763301_300ohm
*******
.subckt 1206_782763480_48ohm 1 2
Rp 1 2 73
Cp 1 2 0.083p
Rs 1 N3 0.005
L1 N3 2 0.084u
.ends 1206_782763480_48ohm
*******
.subckt 1206_782763501_500ohm 1 2
Rp 1 2 550
Cp 1 2 1.179p
Rs 1 N3 0.06
L1 N3 2 1.62u
.ends 1206_782763501_500ohm
*******
.subckt 1206_782763601_600ohm 1 2
Rp 1 2 620
Cp 1 2 1.9p
Rs 1 N3 0.048
L1 N3 2 1.8u
.ends 1206_782763601_600ohm
*******
.subckt 1206_782763621_620ohm 1 2
Rp 1 2 620
Cp 1 2 1.1p
Rs 1 N3 0.1
L1 N3 2 3.2u
.ends 1206_782763621_620ohm
*******
.subckt 1206_782763700_70ohm 1 2
Rp 1 2 100
Cp 1 2 0.145p
Rs 1 N3 0.15
L1 N3 2 0.223u
.ends 1206_782763700_70ohm
*******
.subckt 1206_782763800_80ohm 1 2
Rp 1 2 88
Cp 1 2 0.072p
Rs 1 N3 0.02
L1 N3 2 0.252u
.ends 1206_782763800_80ohm
*******
.subckt 1206_782763820_82ohm 1 2
Rp 1 2 120
Cp 1 2 0.4p
Rs 1 N3 0.025
L1 N3 2 0.275u
.ends 1206_782763820_82ohm
*******
.subckt 1806_782963201_1000ohm 1 2
Rp 1 2 1.273
Cp 1 2 1.049p
Rs 1 N3 0.09
L1 N3 2 0.005396u
.ends 1806_782963201_1000ohm
*******
.subckt 1806_782963560_56ohm 1 2
Rp 1 2 74.5
Cp 1 2 0.102p
Rs 1 N3 0.008
L1 N3 2 0.21u
.ends 1806_782963560_56ohm
*******
.subckt 1806_782963600_60ohm 1 2
Rp 1 2 79.2262562115367
Cp 1 2 72.6079064201p
Rs 1 N3 0.01
L1 N3 2 0.232761224934067u
.ends 1806_782963600_60ohm
*******
.subckt 1806_782963610_60ohm 1 2
Rp 1 2 111
Cp 1 2 0.034p
Rs 1 N3 0.008
L1 N3 2 0.148u
.ends 1806_782963610_60ohm
*******
.subckt 1806_782963800_80ohm 1 2
Rp 1 2 80
Cp 1 2 0.04p
Rs 1 N3 0.04
L1 N3 2 0.3u
.ends 1806_782963800_80ohm
*******
.subckt 1806_782963820_82ohm 1 2
Rp 1 2 87.1
Cp 1 2 0.127p
Rs 1 N3 0.02
L1 N3 2 0.213u
.ends 1806_782963820_82ohm
*******
.subckt 1806_782963851_850ohm 1 2
Rp 1 2 1146
Cp 1 2 2.55p
Rs 1 N3 0.1
L1 N3 2 3.541u
.ends 1806_782963851_850ohm
*******
.subckt 1812_782965121_120ohm 1 2
Rp 1 2 152
Cp 1 2 0.36p
Rs 1 N3 0.04
L1 N3 2 0.482u
.ends 1812_782965121_120ohm
*******
.subckt 1812_782965601_600ohm 1 2
Rp 1 2 981
Cp 1 2 4.9p
Rs 1 N3 0.04
L1 N3 2 1.116u
.ends 1812_782965601_600ohm
*******
.subckt 1812_782965700_70ohm 1 2
Rp 1 2 100
Cp 1 2 0.101p
Rs 1 N3 0.008
L1 N3 2 0.284u
.ends 1812_782965700_70ohm
*******
.subckt 1812_782965781_780ohm 1 2
Rp 1 2 1616
Cp 1 2 3.6p
Rs 1 N3 0.04
L1 N3 2 1.4u
.ends 1812_782965781_780ohm
*******
