**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Optocoupler Phototransistor
* Matchcode:              WL-OCPT
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
********************************************************
***********************Series_10x***********************
********************************************************
***********************
.SUBCKT Series_10x_140105146000 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.44307E+01*PWR(V(T),(0.11596E+01+0.27749E+01*V(T)))-.76712E+00*V(T))/100,
+ (0.82049E-02*(PWR(0.98748E+00,(1/V(T))))*PWR(V(T),-.30962E+00)+0.10511E+00*V(T))/97)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=89.506E-18
+ N=1.4695
+ RS=1.1278
+ IKF=18.225E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=100 NF=1.1 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_10x_140106146000 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.44307E+01*PWR(V(T),(0.11596E+01+0.27749E+01*V(T)))-.76712E+00*V(T))/100,
+ (0.82049E-02*(PWR(0.98748E+00,(1/V(T))))*PWR(V(T),-.30962E+00)+0.10511E+00*V(T))/97)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=89.506E-18
+ N=1.4695
+ RS=1.1278
+ IKF=18.225E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=120 NF=1.1 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_10x_140107146000 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.44307E+01*PWR(V(T),(0.11596E+01+0.27749E+01*V(T)))-.76712E+00*V(T))/100,
+ (0.82049E-02*(PWR(0.98748E+00,(1/V(T))))*PWR(V(T),-.30962E+00)+0.10511E+00*V(T))/97)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=89.506E-18
+ N=1.4695
+ RS=1.1278
+ IKF=18.225E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=200 NF=1.1 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_10x_140108146000 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.44307E+01*PWR(V(T),(0.11596E+01+0.27749E+01*V(T)))-.76712E+00*V(T))/100,
+ (0.82049E-02*(PWR(0.98748E+00,(1/V(T))))*PWR(V(T),-.30962E+00)+0.10511E+00*V(T))/97)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=89.506E-18
+ N=1.4695
+ RS=1.1278
+ IKF=18.225E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=200 NF=1.1 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_10x_140109146000 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.44307E+01*PWR(V(T),(0.11596E+01+0.27749E+01*V(T)))-.76712E+00*V(T))/100,
+ (0.82049E-02*(PWR(0.98748E+00,(1/V(T))))*PWR(V(T),-.30962E+00)+0.10511E+00*V(T))/97)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=89.506E-18
+ N=1.4695
+ RS=1.1278
+ IKF=18.225E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=300 NF=1.1 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_10x_140100146000 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.44307E+01*PWR(V(T),(0.11596E+01+0.27749E+01*V(T)))-.76712E+00*V(T))/100,
+ (0.82049E-02*(PWR(0.98748E+00,(1/V(T))))*PWR(V(T),-.30962E+00)+0.10511E+00*V(T))/97)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=89.506E-18
+ N=1.4695
+ RS=1.1278
+ IKF=18.225E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=450 NF=1.1 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
********************************************************
***********************Series_354***********************
********************************************************
***********************
.SUBCKT Series_354_140354245100 A K C E 
D1 A D LED
VH D K 0 
Hd R 0 VH 1
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.02,
+ ((0.43970E+01-.21363E-04*PWR(V(T),-.12107E+01))/(0.18799E+02+PWR(V(T),-.12107E+01)))/100,
+ (1/(0.87599E+02*PWR((V(T)+0.11261E-01),2)+0.63063E+01)+0.31648E-01*Ln(V(T)))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=31.851E-18
+ N=1.4226
+ RS=.71497
+ IKF=11.194E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=150 NF=1.14 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=65 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_354_140354245000 A K C E 
D1 A D LED
VH D K 0 
Hd R 0 VH 1
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.02,
+ ((0.43970E+01-.21363E-04*PWR(V(T),-.12107E+01))/(0.18799E+02+PWR(V(T),-.12107E+01)))/100,
+ (1/(0.87599E+02*PWR((V(T)+0.11261E-01),2)+0.63063E+01)+0.31648E-01*Ln(V(T)))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=31.851E-18
+ N=1.4226
+ RS=.71497
+ IKF=11.194E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=150 NF=1.14 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=65 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
********************************************************
***********************Series_356***********************
********************************************************
***********************
.SUBCKT Series_356_140356145000 A K C E 
D1 A D LED
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=100 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_356_140356145100 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=120 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_356_140356145200 A K C E 
D1 A D LED
VH D K 0
Hd R 0 VH 1
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=200 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_356_140356145300 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=300 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_356_140356145400 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=450 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
********************************************************
***********************Series_357***********************
********************************************************
***********************
.SUBCKT Series_357_140357145000 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=350 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_357_140357145100 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=120 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_357_140357145200 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=200 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_357_140357145300 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=300 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_357_140357145400 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.025,
+ (0.87984E+01*PWR(V(T),(0.13437E+01+0.38089E+01*V(T)))-.28829E+00*V(T))/100,
+ (0.19311E+05*PWR(V(T),(0.29342E+01+0.29886E+02*V(T)))+0.46089E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=6.9809E-15
+ N=1.6332
+ RS=1.8224
+ IKF=.10986
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=450 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
********************************************************
***********************Series_814***********************
********************************************************
***********************
.SUBCKT Series_814_14081424x1x0 A K C E 
D1 A D LED
VH D K 0 
Hd R 0 VH 1
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.015,
+ (0.76070E+01*PWR(V(T),(0.12094E+01+0.26644E+01*V(T)))-.76178E+00*V(T))/100,
+ (0.10247E+04*PWR(V(T),(0.21850E+01+0.26273E+02*V(T)))+0.53977E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=87.786E-18
+ N=1.4594
+ RS=1.1118
+ IKF=160.02
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=100 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=65 IKF=1 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_814_14081424x0x0 A K C E 
D1 A D LED
VH D K 0 
Hd R 0 VH 1
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.015,
+ (0.76070E+01*PWR(V(T),(0.12094E+01+0.26644E+01*V(T)))-.76178E+00*V(T))/100,
+ (0.10247E+04*PWR(V(T),(0.21850E+01+0.26273E+02*V(T)))+0.53977E+00*V(T))/99)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=87.786E-18
+ N=1.4594
+ RS=1.1118
+ IKF=160.02
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=150 NF=1.145 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=65 IKF=1 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
********************************************************
***********************Series_816***********************
********************************************************
***********************
.SUBCKT Series_816_14081614x0x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=350 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_816_14081614x1x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=120 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_816_14081614x2x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=200 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_816_14081614x3x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=300 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_816_14081614x4x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=450 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
********************************************************
***********************Series_817***********************
********************************************************
***********************
.SUBCKT Series_817_14081714x0x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=350 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_817_14081714x1x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=120 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_817_14081714x2x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=200 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_817_14081714x3x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=300 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_817_14081714x4x0 A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector 

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.49207E+01*PWR(V(T),(0.11893E+01+0.38933E+01*V(T)))-.62825E+00*V(T))/100,
+ (-.23752E-01*EXP(-.11157E+03*V(T))+0.17792E-01*EXP(0.30610E+01*V(T)))/96.5)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=1.1516E-15
+ N=1.6015
+ RS=2.0027
+ IKF=19.785E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=450 NF=1.13 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=0.5 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_827_14082718xxx A K C E A1 K1 C1 E1 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.01,
+ (0.75567E+01*PWR(V(T),(0.12975E+01+0.48156E+01*V(T)))-.37487E+00*V(T) )/100,
+ (0.19358E-01*EXP((PWR((Ln(V(T))+.34026E+01),2))/-.18146E+01)+0.29107E+00*V(T))/100)}
+ (0,0.0000000001) (10,10)

D2 A1 D1 LED	
VH1 D1 K1 0 
Hd1 R1 0 VH1 1	
Rd1 R1 T1 10k
Cd1 T1 0 0.02n
Rg1 B1 0 4G
Q2 C1 B1 E1 Detector

G2 C1 B1 TABLE
+ {if(V(T1)<0.01,
+ (0.75567E+01*PWR(V(T1),(0.12975E+01+0.48156E+01*V(T1)))-.37487E+00*V(T1) )/100,
+ (0.19358E-01*EXP((PWR((Ln(V(T1))+.34026E+01),2))/-.18146E+01)+0.29107E+00*V(T1))/100)}
+ (0,0.0000000001) (10,10)

.model LED D 
+ IS=209.97E-18
+ N=1.5072
+ RS=1.1904
+ IKF=.30047
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9
.model Detector NPN IS=3.64P BF=625 NF=1.3 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=10 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************