**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Infrared TOP LED Waterclear
* Matchcode:              WL-SITW
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-03-02
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 3528_15414185BA210 1 2
D1 1 2 led
.MODEL led D
+ IS=124.66E-21
+ N=1.3198
+ RS=.90718
+ IKF=66.101E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*******
.subckt 3528_15414194BA210 1 2
D1 1 2 led
.MODEL led D
+ IS=1.3840E-15
+ N=1.6688
+ RS=1.6640
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*******
.subckt 3528_15414185A3011 1 2
D1 1 2 led
.MODEL led D
+ IS=3.1747E-18
+ N=1.4492
+ RS=1.3797
+ IKF=30.726E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*******
.subckt 3528_15414185A6011 1 2
D1 1 2 led
.MODEL led D
+ IS=3.3666E-18
+ N=1.4497
+ RS=1.8735
+ IKF=13.191E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*******
.subckt 3528_15414185AA211 1 2
D1 1 2 led
.MODEL led D
+ IS=2.4731E-18
+ N=1.4363
+ RS=1.5712
+ IKF=27.574E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*******
.subckt 3528_15414194A3011 1 2
D1 1 2 led
.MODEL led D
+ IS=8.9658E-18
+ N=1.3401
+ RS=1.1998
+ IKF=14.406E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*******
.subckt 3528_15414194A6011 1 2
D1 1 2 led
.MODEL led D
+ IS=10.205E-18
+ N=1.3470
+ RS=1.1736
+ IKF=14.608E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*******
.subckt 3528_15414194AA211 1 2
D1 1 2 led
.MODEL led D
+ IS=12.486E-18
+ N=1.3538
+ RS=.74728
+ IKF=53.166E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=100.00E-6
.ends
*******

































