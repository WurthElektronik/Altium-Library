**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Ceramic Common Mode Filter
* Matchcode:              WE-CCMF 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt WE-CCMF_748020024 1 2 3 4
Vam1 1 n2 dc 0
Rport1 n2 0 50
Vam2 2 n4 dc 0
Rport2 n4 0 50
Vam3 3 n6 dc 0
Rport3 n6 0 50
Vam4 4 n8 dc 0
Rport4 n8 0 50

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1
Fi3 0 ni3 Vam3 50
Gi3 0 ni3 3 0 1
Rt3 ni3 0 1
Fi4 0 ni4 Vam4 50
Gi4 0 ni4 4 0 1
Rt4 ni4 0 1

Ca1 ns1 0 1e-012
Ca2 ns2 0 1e-012
Ra1 ns1 0 147.219400304
Ra2 ns2 0 147.219400304
Ga1 ns1 0 ns2 0 -0.00204136883855
Ga2 ns2 0 ns1 0 0.00204136883855
Ca3 ns3 0 1e-012
Ca4 ns4 0 1e-012
Ra3 ns3 0 229.546477593
Ra4 ns4 0 229.546477593
Ga3 ns3 0 ns4 0 -0.00836983773395
Ga4 ns4 0 ns3 0 0.00836983773395
Ca5 ns5 0 1e-012
Ca6 ns6 0 1e-012
Ra5 ns5 0 145.303135369
Ra6 ns6 0 145.303135369
Ga5 ns5 0 ns6 0 -0.0221791727372
Ga6 ns6 0 ns5 0 0.0221791727372
Ca7 ns7 0 1e-012
Ca8 ns8 0 1e-012
Ra7 ns7 0 125.51202363
Ra8 ns8 0 125.51202363
Ga7 ns7 0 ns8 0 -0.0390361561464
Ga8 ns8 0 ns7 0 0.0390361561464
Ca9 ns9 0 1e-012
Ca10 ns10 0 1e-012
Ra9 ns9 0 1099.82097604
Ra10 ns10 0 1099.82097604
Ga9 ns9 0 ns10 0 -0.0431338846321
Ga10 ns10 0 ns9 0 0.0431338846321
Ca11 ns11 0 1e-012
Ca12 ns12 0 1e-012
Ra11 ns11 0 89.6349355902
Ra12 ns12 0 89.6349355902
Ga11 ns11 0 ns12 0 -0.0527305240232
Ga12 ns12 0 ns11 0 0.0527305240232
Ca13 ns13 0 1e-012
Ca14 ns14 0 1e-012
Ra13 ns13 0 116.544388093
Ra14 ns14 0 116.544388093
Ga13 ns13 0 ns14 0 -0.0596819754204
Ga14 ns14 0 ns13 0 0.0596819754204
Ca15 ns15 0 1e-012
Ca16 ns16 0 1e-012
Ra15 ns15 0 157.874603033
Ra16 ns16 0 157.874603033
Ga15 ns15 0 ns16 0 -0.070138824588
Ga16 ns16 0 ns15 0 0.070138824588
Ca17 ns17 0 1e-012
Ca18 ns18 0 1e-012
Ra17 ns17 0 185.317195465
Ra18 ns18 0 185.317195465
Ga17 ns17 0 ns18 0 -0.073707531923
Ga18 ns18 0 ns17 0 0.073707531923
Ca19 ns19 0 1e-012
Ca20 ns20 0 1e-012
Ra19 ns19 0 138.938682675
Ra20 ns20 0 138.938682675
Ga19 ns19 0 ns20 0 -0.0818972981799
Ga20 ns20 0 ns19 0 0.0818972981799
Ca21 ns21 0 1e-012
Ca22 ns22 0 1e-012
Ra21 ns21 0 176.387891511
Ra22 ns22 0 176.387891511
Ga21 ns21 0 ns22 0 -0.0916634820428
Ga22 ns22 0 ns21 0 0.0916634820428
Ca23 ns23 0 1e-012
Ca24 ns24 0 1e-012
Ra23 ns23 0 147.219400304
Ra24 ns24 0 147.219400304
Ga23 ns23 0 ns24 0 -0.00204136883855
Ga24 ns24 0 ns23 0 0.00204136883855
Ca25 ns25 0 1e-012
Ca26 ns26 0 1e-012
Ra25 ns25 0 229.546477593
Ra26 ns26 0 229.546477593
Ga25 ns25 0 ns26 0 -0.00836983773395
Ga26 ns26 0 ns25 0 0.00836983773395
Ca27 ns27 0 1e-012
Ca28 ns28 0 1e-012
Ra27 ns27 0 145.303135369
Ra28 ns28 0 145.303135369
Ga27 ns27 0 ns28 0 -0.0221791727372
Ga28 ns28 0 ns27 0 0.0221791727372
Ca29 ns29 0 1e-012
Ca30 ns30 0 1e-012
Ra29 ns29 0 125.51202363
Ra30 ns30 0 125.51202363
Ga29 ns29 0 ns30 0 -0.0390361561464
Ga30 ns30 0 ns29 0 0.0390361561464
Ca31 ns31 0 1e-012
Ca32 ns32 0 1e-012
Ra31 ns31 0 1099.82097604
Ra32 ns32 0 1099.82097604
Ga31 ns31 0 ns32 0 -0.0431338846321
Ga32 ns32 0 ns31 0 0.0431338846321
Ca33 ns33 0 1e-012
Ca34 ns34 0 1e-012
Ra33 ns33 0 89.6349355902
Ra34 ns34 0 89.6349355902
Ga33 ns33 0 ns34 0 -0.0527305240232
Ga34 ns34 0 ns33 0 0.0527305240232
Ca35 ns35 0 1e-012
Ca36 ns36 0 1e-012
Ra35 ns35 0 116.544388093
Ra36 ns36 0 116.544388093
Ga35 ns35 0 ns36 0 -0.0596819754204
Ga36 ns36 0 ns35 0 0.0596819754204
Ca37 ns37 0 1e-012
Ca38 ns38 0 1e-012
Ra37 ns37 0 157.874603033
Ra38 ns38 0 157.874603033
Ga37 ns37 0 ns38 0 -0.070138824588
Ga38 ns38 0 ns37 0 0.070138824588
Ca39 ns39 0 1e-012
Ca40 ns40 0 1e-012
Ra39 ns39 0 185.317195465
Ra40 ns40 0 185.317195465
Ga39 ns39 0 ns40 0 -0.073707531923
Ga40 ns40 0 ns39 0 0.073707531923
Ca41 ns41 0 1e-012
Ca42 ns42 0 1e-012
Ra41 ns41 0 138.938682675
Ra42 ns42 0 138.938682675
Ga41 ns41 0 ns42 0 -0.0818972981799
Ga42 ns42 0 ns41 0 0.0818972981799
Ca43 ns43 0 1e-012
Ca44 ns44 0 1e-012
Ra43 ns43 0 176.387891511
Ra44 ns44 0 176.387891511
Ga43 ns43 0 ns44 0 -0.0916634820428
Ga44 ns44 0 ns43 0 0.0916634820428
Ca45 ns45 0 1e-012
Ca46 ns46 0 1e-012
Ra45 ns45 0 147.219400304
Ra46 ns46 0 147.219400304
Ga45 ns45 0 ns46 0 -0.00204136883855
Ga46 ns46 0 ns45 0 0.00204136883855
Ca47 ns47 0 1e-012
Ca48 ns48 0 1e-012
Ra47 ns47 0 229.546477593
Ra48 ns48 0 229.546477593
Ga47 ns47 0 ns48 0 -0.00836983773395
Ga48 ns48 0 ns47 0 0.00836983773395
Ca49 ns49 0 1e-012
Ca50 ns50 0 1e-012
Ra49 ns49 0 145.303135369
Ra50 ns50 0 145.303135369
Ga49 ns49 0 ns50 0 -0.0221791727372
Ga50 ns50 0 ns49 0 0.0221791727372
Ca51 ns51 0 1e-012
Ca52 ns52 0 1e-012
Ra51 ns51 0 125.51202363
Ra52 ns52 0 125.51202363
Ga51 ns51 0 ns52 0 -0.0390361561464
Ga52 ns52 0 ns51 0 0.0390361561464
Ca53 ns53 0 1e-012
Ca54 ns54 0 1e-012
Ra53 ns53 0 1099.82097604
Ra54 ns54 0 1099.82097604
Ga53 ns53 0 ns54 0 -0.0431338846321
Ga54 ns54 0 ns53 0 0.0431338846321
Ca55 ns55 0 1e-012
Ca56 ns56 0 1e-012
Ra55 ns55 0 89.6349355902
Ra56 ns56 0 89.6349355902
Ga55 ns55 0 ns56 0 -0.0527305240232
Ga56 ns56 0 ns55 0 0.0527305240232
Ca57 ns57 0 1e-012
Ca58 ns58 0 1e-012
Ra57 ns57 0 116.544388093
Ra58 ns58 0 116.544388093
Ga57 ns57 0 ns58 0 -0.0596819754204
Ga58 ns58 0 ns57 0 0.0596819754204
Ca59 ns59 0 1e-012
Ca60 ns60 0 1e-012
Ra59 ns59 0 157.874603033
Ra60 ns60 0 157.874603033
Ga59 ns59 0 ns60 0 -0.070138824588
Ga60 ns60 0 ns59 0 0.070138824588
Ca61 ns61 0 1e-012
Ca62 ns62 0 1e-012
Ra61 ns61 0 185.317195465
Ra62 ns62 0 185.317195465
Ga61 ns61 0 ns62 0 -0.073707531923
Ga62 ns62 0 ns61 0 0.073707531923
Ca63 ns63 0 1e-012
Ca64 ns64 0 1e-012
Ra63 ns63 0 138.938682675
Ra64 ns64 0 138.938682675
Ga63 ns63 0 ns64 0 -0.0818972981799
Ga64 ns64 0 ns63 0 0.0818972981799
Ca65 ns65 0 1e-012
Ca66 ns66 0 1e-012
Ra65 ns65 0 176.387891511
Ra66 ns66 0 176.387891511
Ga65 ns65 0 ns66 0 -0.0916634820428
Ga66 ns66 0 ns65 0 0.0916634820428
Ca67 ns67 0 1e-012
Ca68 ns68 0 1e-012
Ra67 ns67 0 147.219400304
Ra68 ns68 0 147.219400304
Ga67 ns67 0 ns68 0 -0.00204136883855
Ga68 ns68 0 ns67 0 0.00204136883855
Ca69 ns69 0 1e-012
Ca70 ns70 0 1e-012
Ra69 ns69 0 229.546477593
Ra70 ns70 0 229.546477593
Ga69 ns69 0 ns70 0 -0.00836983773395
Ga70 ns70 0 ns69 0 0.00836983773395
Ca71 ns71 0 1e-012
Ca72 ns72 0 1e-012
Ra71 ns71 0 145.303135369
Ra72 ns72 0 145.303135369
Ga71 ns71 0 ns72 0 -0.0221791727372
Ga72 ns72 0 ns71 0 0.0221791727372
Ca73 ns73 0 1e-012
Ca74 ns74 0 1e-012
Ra73 ns73 0 125.51202363
Ra74 ns74 0 125.51202363
Ga73 ns73 0 ns74 0 -0.0390361561464
Ga74 ns74 0 ns73 0 0.0390361561464
Ca75 ns75 0 1e-012
Ca76 ns76 0 1e-012
Ra75 ns75 0 1099.82097604
Ra76 ns76 0 1099.82097604
Ga75 ns75 0 ns76 0 -0.0431338846321
Ga76 ns76 0 ns75 0 0.0431338846321
Ca77 ns77 0 1e-012
Ca78 ns78 0 1e-012
Ra77 ns77 0 89.6349355902
Ra78 ns78 0 89.6349355902
Ga77 ns77 0 ns78 0 -0.0527305240232
Ga78 ns78 0 ns77 0 0.0527305240232
Ca79 ns79 0 1e-012
Ca80 ns80 0 1e-012
Ra79 ns79 0 116.544388093
Ra80 ns80 0 116.544388093
Ga79 ns79 0 ns80 0 -0.0596819754204
Ga80 ns80 0 ns79 0 0.0596819754204
Ca81 ns81 0 1e-012
Ca82 ns82 0 1e-012
Ra81 ns81 0 157.874603033
Ra82 ns82 0 157.874603033
Ga81 ns81 0 ns82 0 -0.070138824588
Ga82 ns82 0 ns81 0 0.070138824588
Ca83 ns83 0 1e-012
Ca84 ns84 0 1e-012
Ra83 ns83 0 185.317195465
Ra84 ns84 0 185.317195465
Ga83 ns83 0 ns84 0 -0.073707531923
Ga84 ns84 0 ns83 0 0.073707531923
Ca85 ns85 0 1e-012
Ca86 ns86 0 1e-012
Ra85 ns85 0 138.938682675
Ra86 ns86 0 138.938682675
Ga85 ns85 0 ns86 0 -0.0818972981799
Ga86 ns86 0 ns85 0 0.0818972981799
Ca87 ns87 0 1e-012
Ca88 ns88 0 1e-012
Ra87 ns87 0 176.387891511
Ra88 ns88 0 176.387891511
Ga87 ns87 0 ns88 0 -0.0916634820428
Ga88 ns88 0 ns87 0 0.0916634820428

Gb1_1 ns1 0 ni1 0 0.00740607376079
Gb3_1 ns3 0 ni1 0 0.0106373084965
Gb5_1 ns5 0 ni1 0 0.0243146978621
Gb7_1 ns7 0 ni1 0 0.0406623124611
Gb9_1 ns9 0 ni1 0 0.0431530508946
Gb11_1 ns11 0 ni1 0 0.0550909114427
Gb13_1 ns13 0 ni1 0 0.060915574619
Gb15_1 ns15 0 ni1 0 0.0707108521743
Gb17_1 ns17 0 ni1 0 0.0741025861314
Gb19_1 ns19 0 ni1 0 0.082529832467
Gb21_1 ns21 0 ni1 0 0.0920141258003
Gb23_2 ns23 0 ni2 0 0.00740607376079
Gb25_2 ns25 0 ni2 0 0.0106373084965
Gb27_2 ns27 0 ni2 0 0.0243146978621
Gb29_2 ns29 0 ni2 0 0.0406623124611
Gb31_2 ns31 0 ni2 0 0.0431530508946
Gb33_2 ns33 0 ni2 0 0.0550909114427
Gb35_2 ns35 0 ni2 0 0.060915574619
Gb37_2 ns37 0 ni2 0 0.0707108521743
Gb39_2 ns39 0 ni2 0 0.0741025861314
Gb41_2 ns41 0 ni2 0 0.082529832467
Gb43_2 ns43 0 ni2 0 0.0920141258003
Gb45_3 ns45 0 ni3 0 0.00740607376079
Gb47_3 ns47 0 ni3 0 0.0106373084965
Gb49_3 ns49 0 ni3 0 0.0243146978621
Gb51_3 ns51 0 ni3 0 0.0406623124611
Gb53_3 ns53 0 ni3 0 0.0431530508946
Gb55_3 ns55 0 ni3 0 0.0550909114427
Gb57_3 ns57 0 ni3 0 0.060915574619
Gb59_3 ns59 0 ni3 0 0.0707108521743
Gb61_3 ns61 0 ni3 0 0.0741025861314
Gb63_3 ns63 0 ni3 0 0.082529832467
Gb65_3 ns65 0 ni3 0 0.0920141258003
Gb67_4 ns67 0 ni4 0 0.00740607376079
Gb69_4 ns69 0 ni4 0 0.0106373084965
Gb71_4 ns71 0 ni4 0 0.0243146978621
Gb73_4 ns73 0 ni4 0 0.0406623124611
Gb75_4 ns75 0 ni4 0 0.0431530508946
Gb77_4 ns77 0 ni4 0 0.0550909114427
Gb79_4 ns79 0 ni4 0 0.060915574619
Gb81_4 ns81 0 ni4 0 0.0707108521743
Gb83_4 ns83 0 ni4 0 0.0741025861314
Gb85_4 ns85 0 ni4 0 0.082529832467
Gb87_4 ns87 0 ni4 0 0.0920141258003

Gc1_1 0 n2 ns1 0 -0.0481253057691
Gc1_2 0 n2 ns2 0 -0.0596402932528
Gc1_3 0 n2 ns3 0 0.00752736067566
Gc1_4 0 n2 ns4 0 -0.0074084118514
Gc1_5 0 n2 ns5 0 -0.0113650667706
Gc1_6 0 n2 ns6 0 -0.00394231073944
Gc1_7 0 n2 ns7 0 -0.00229949444909
Gc1_8 0 n2 ns8 0 -0.00131757923003
Gc1_9 0 n2 ns9 0 -9.84363258406e-005
Gc1_10 0 n2 ns10 0 2.7523488714e-005
Gc1_11 0 n2 ns11 0 -0.00627006930415
Gc1_12 0 n2 ns12 0 0.00922495737249
Gc1_13 0 n2 ns13 0 -0.0089975603813
Gc1_14 0 n2 ns14 0 -0.00893855898535
Gc1_15 0 n2 ns15 0 0.00152653865379
Gc1_16 0 n2 ns16 0 -0.000819302602467
Gc1_17 0 n2 ns17 0 -0.00167074451981
Gc1_18 0 n2 ns18 0 -0.00285085644892
Gc1_19 0 n2 ns19 0 6.67231332448e-006
Gc1_20 0 n2 ns20 0 -0.00156451109989
Gc1_21 0 n2 ns21 0 -0.000301226398416
Gc1_22 0 n2 ns22 0 -0.000473910797718
Gc1_23 0 n2 ns23 0 0.013609690519
Gc1_24 0 n2 ns24 0 0.00463953759832
Gc1_25 0 n2 ns25 0 0.00952180445444
Gc1_26 0 n2 ns26 0 0.00394434388338
Gc1_27 0 n2 ns27 0 0.00133507073509
Gc1_28 0 n2 ns28 0 -0.000225883397833
Gc1_29 0 n2 ns29 0 0.00383317429164
Gc1_30 0 n2 ns30 0 0.00322223383552
Gc1_31 0 n2 ns31 0 -4.22222627333e-005
Gc1_32 0 n2 ns32 0 3.47366293412e-006
Gc1_33 0 n2 ns33 0 -0.000728275696648
Gc1_34 0 n2 ns34 0 -0.00660155748911
Gc1_35 0 n2 ns35 0 0.00465981660769
Gc1_36 0 n2 ns36 0 0.00329438818996
Gc1_37 0 n2 ns37 0 0.00646348929953
Gc1_38 0 n2 ns38 0 0.00218243712696
Gc1_39 0 n2 ns39 0 -0.00388427613035
Gc1_40 0 n2 ns40 0 0.00244625762359
Gc1_41 0 n2 ns41 0 -0.000141670783265
Gc1_42 0 n2 ns42 0 0.000739811499601
Gc1_43 0 n2 ns43 0 -0.000837939513942
Gc1_44 0 n2 ns44 0 0.00114455422267
Gc1_45 0 n2 ns45 0 -0.00196742747959
Gc1_46 0 n2 ns46 0 0.0128610310469
Gc1_47 0 n2 ns47 0 0.00564334343304
Gc1_48 0 n2 ns48 0 0.00915868592321
Gc1_49 0 n2 ns49 0 0.0102118091476
Gc1_50 0 n2 ns50 0 0.000634081855902
Gc1_51 0 n2 ns51 0 -0.00167158094478
Gc1_52 0 n2 ns52 0 -0.00314987499513
Gc1_53 0 n2 ns53 0 6.45753418973e-005
Gc1_54 0 n2 ns54 0 -2.17649889982e-005
Gc1_55 0 n2 ns55 0 0.001506477089
Gc1_56 0 n2 ns56 0 0.00215066248408
Gc1_57 0 n2 ns57 0 0.00421891676213
Gc1_58 0 n2 ns58 0 0.00492338744356
Gc1_59 0 n2 ns59 0 -7.6953297705e-005
Gc1_60 0 n2 ns60 0 0.00165850467171
Gc1_61 0 n2 ns61 0 -0.00103416013108
Gc1_62 0 n2 ns62 0 -0.00127534396565
Gc1_63 0 n2 ns63 0 -0.00151261811196
Gc1_64 0 n2 ns64 0 0.00123632577124
Gc1_65 0 n2 ns65 0 -0.000312330103352
Gc1_66 0 n2 ns66 0 0.000891567867762
Gc1_67 0 n2 ns67 0 0.0143265553778
Gc1_68 0 n2 ns68 0 0.00672122682366
Gc1_69 0 n2 ns69 0 0.00872257514111
Gc1_70 0 n2 ns70 0 0.00470395130504
Gc1_71 0 n2 ns71 0 0.000660357112417
Gc1_72 0 n2 ns72 0 -0.000293258802625
Gc1_73 0 n2 ns73 0 0.00205256177245
Gc1_74 0 n2 ns74 0 0.00278156027639
Gc1_75 0 n2 ns75 0 5.73082404113e-005
Gc1_76 0 n2 ns76 0 -1.02757589666e-005
Gc1_77 0 n2 ns77 0 0.00465054778114
Gc1_78 0 n2 ns78 0 0.00280033870859
Gc1_79 0 n2 ns79 0 -0.00159970462656
Gc1_80 0 n2 ns80 0 0.000268846819924
Gc1_81 0 n2 ns81 0 0.000595336651121
Gc1_82 0 n2 ns82 0 0.00281957549478
Gc1_83 0 n2 ns83 0 -0.000911173414912
Gc1_84 0 n2 ns84 0 5.67533191682e-005
Gc1_85 0 n2 ns85 0 -0.000874289752461
Gc1_86 0 n2 ns86 0 0.000760347075436
Gc1_87 0 n2 ns87 0 0.000637887123607
Gc1_88 0 n2 ns88 0 -0.000442499808627
Gd1_1 0 n2 ni1 0 -0.0150756254366
Gd1_2 0 n2 ni2 0 0.00896002734602
Gd1_3 0 n2 ni3 0 0.00416062326128
Gd1_4 0 n2 ni4 0 0.00473339222916
Gc2_1 0 n4 ns1 0 0.0136664032411
Gc2_2 0 n4 ns2 0 0.00467809277143
Gc2_3 0 n4 ns3 0 0.00953608135482
Gc2_4 0 n4 ns4 0 0.00395720732544
Gc2_5 0 n4 ns5 0 0.00134689592354
Gc2_6 0 n4 ns6 0 -0.000229067747563
Gc2_7 0 n4 ns7 0 0.00385631604085
Gc2_8 0 n4 ns8 0 0.00321956752141
Gc2_9 0 n4 ns9 0 -4.21916697085e-005
Gc2_10 0 n4 ns10 0 3.72864248341e-006
Gc2_11 0 n4 ns11 0 -0.000690076685458
Gc2_12 0 n4 ns12 0 -0.00657639840027
Gc2_13 0 n4 ns13 0 0.00463850952013
Gc2_14 0 n4 ns14 0 0.00331329739265
Gc2_15 0 n4 ns15 0 0.00646727090811
Gc2_16 0 n4 ns16 0 0.00218812473025
Gc2_17 0 n4 ns17 0 -0.0038947492028
Gc2_18 0 n4 ns18 0 0.00244900311738
Gc2_19 0 n4 ns19 0 -0.000147966106615
Gc2_20 0 n4 ns20 0 0.000736605599077
Gc2_21 0 n4 ns21 0 -0.000840400081286
Gc2_22 0 n4 ns22 0 0.00114493141547
Gc2_23 0 n4 ns23 0 -0.0106144384664
Gc2_24 0 n4 ns24 0 -0.00818390841432
Gc2_25 0 n4 ns25 0 0.00752247639657
Gc2_26 0 n4 ns26 0 0.00582850491057
Gc2_27 0 n4 ns27 0 -0.012677754283
Gc2_28 0 n4 ns28 0 0.000924385148274
Gc2_29 0 n4 ns29 0 -0.00318885717456
Gc2_30 0 n4 ns30 0 -0.00293100446684
Gc2_31 0 n4 ns31 0 -5.45538625535e-005
Gc2_32 0 n4 ns32 0 2.30789956037e-005
Gc2_33 0 n4 ns33 0 0.000276674062965
Gc2_34 0 n4 ns34 0 0.0042806831622
Gc2_35 0 n4 ns35 0 -0.00669253260903
Gc2_36 0 n4 ns36 0 -0.00387190752321
Gc2_37 0 n4 ns37 0 0.00506361867839
Gc2_38 0 n4 ns38 0 0.00293341899973
Gc2_39 0 n4 ns39 0 -0.00439437950939
Gc2_40 0 n4 ns40 0 -0.00200416960091
Gc2_41 0 n4 ns41 0 -0.00215317507371
Gc2_42 0 n4 ns42 0 -0.000696027398857
Gc2_43 0 n4 ns43 0 -0.000360373647221
Gc2_44 0 n4 ns44 0 -0.000282162140293
Gc2_45 0 n4 ns45 0 0.0157058424033
Gc2_46 0 n4 ns46 0 0.00723893927849
Gc2_47 0 n4 ns47 0 0.00939294286136
Gc2_48 0 n4 ns48 0 0.00476430115531
Gc2_49 0 n4 ns49 0 0.00137748257137
Gc2_50 0 n4 ns50 0 -0.000136708565665
Gc2_51 0 n4 ns51 0 0.00195862100593
Gc2_52 0 n4 ns52 0 0.00233201611015
Gc2_53 0 n4 ns53 0 5.89774606979e-005
Gc2_54 0 n4 ns54 0 -5.38910114983e-006
Gc2_55 0 n4 ns55 0 0.00785317924429
Gc2_56 0 n4 ns56 0 0.00137141626393
Gc2_57 0 n4 ns57 0 -0.00183781862018
Gc2_58 0 n4 ns58 0 0.00327684902246
Gc2_59 0 n4 ns59 0 -0.000817102213878
Gc2_60 0 n4 ns60 0 0.002484548931
Gc2_61 0 n4 ns61 0 -0.000599552149635
Gc2_62 0 n4 ns62 0 -0.000101247422086
Gc2_63 0 n4 ns63 0 -0.000622289866519
Gc2_64 0 n4 ns64 0 0.00089867139158
Gc2_65 0 n4 ns65 0 0.000571158747285
Gc2_66 0 n4 ns66 0 -1.58124096369e-006
Gc2_67 0 n4 ns67 0 -0.00771495995578
Gc2_68 0 n4 ns68 0 0.00709576434391
Gc2_69 0 n4 ns69 0 0.00570531084256
Gc2_70 0 n4 ns70 0 0.00686680319246
Gc2_71 0 n4 ns71 0 0.00935082636571
Gc2_72 0 n4 ns72 0 -0.00119010986338
Gc2_73 0 n4 ns73 0 -0.00214316252798
Gc2_74 0 n4 ns74 0 -0.00277305168909
Gc2_75 0 n4 ns75 0 5.92832172229e-005
Gc2_76 0 n4 ns76 0 -5.89156078934e-006
Gc2_77 0 n4 ns77 0 0.00182273741779
Gc2_78 0 n4 ns78 0 0.00244972210709
Gc2_79 0 n4 ns79 0 0.00442159791602
Gc2_80 0 n4 ns80 0 0.00347726587611
Gc2_81 0 n4 ns81 0 -0.000863251301323
Gc2_82 0 n4 ns82 0 0.00123163032798
Gc2_83 0 n4 ns83 0 -0.000304664810963
Gc2_84 0 n4 ns84 0 -0.00124519994314
Gc2_85 0 n4 ns85 0 -0.000961311455468
Gc2_86 0 n4 ns86 0 0.0024138910578
Gc2_87 0 n4 ns87 0 -0.000379735007065
Gc2_88 0 n4 ns88 0 0.000645563157363
Gd2_1 0 n4 ni1 0 0.00896780307422
Gd2_2 0 n4 ni2 0 -0.0135138846614
Gd2_3 0 n4 ni3 0 0.0056307464846
Gd2_4 0 n4 ni4 0 0.00340028157587
Gc3_1 0 n6 ns1 0 -0.00186962065562
Gc3_2 0 n6 ns2 0 0.012995147315
Gc3_3 0 n6 ns3 0 0.00563645385865
Gc3_4 0 n6 ns4 0 0.00918803373897
Gc3_5 0 n6 ns5 0 0.0102356839252
Gc3_6 0 n6 ns6 0 0.000641346414804
Gc3_7 0 n6 ns7 0 -0.00166394043586
Gc3_8 0 n6 ns8 0 -0.00314135823511
Gc3_9 0 n6 ns9 0 6.48232574069e-005
Gc3_10 0 n6 ns10 0 -2.17537763e-005
Gc3_11 0 n6 ns11 0 0.00151485091789
Gc3_12 0 n6 ns12 0 0.00215932416695
Gc3_13 0 n6 ns13 0 0.00422645633363
Gc3_14 0 n6 ns14 0 0.00495933686252
Gc3_15 0 n6 ns15 0 -0.000102529392153
Gc3_16 0 n6 ns16 0 0.0016750438224
Gc3_17 0 n6 ns17 0 -0.00104015381635
Gc3_18 0 n6 ns18 0 -0.00129399947062
Gc3_19 0 n6 ns19 0 -0.00151729788745
Gc3_20 0 n6 ns20 0 0.00123319887898
Gc3_21 0 n6 ns21 0 -0.000311176068949
Gc3_22 0 n6 ns22 0 0.00089065270453
Gc3_23 0 n6 ns23 0 0.0156113065654
Gc3_24 0 n6 ns24 0 0.00714358931567
Gc3_25 0 n6 ns25 0 0.00939119240311
Gc3_26 0 n6 ns26 0 0.00473753538432
Gc3_27 0 n6 ns27 0 0.00136393937206
Gc3_28 0 n6 ns28 0 -0.000141484188049
Gc3_29 0 n6 ns29 0 0.00194427241002
Gc3_30 0 n6 ns30 0 0.00232775040735
Gc3_31 0 n6 ns31 0 5.90818106547e-005
Gc3_32 0 n6 ns32 0 -5.34097690405e-006
Gc3_33 0 n6 ns33 0 0.00784126007089
Gc3_34 0 n6 ns34 0 0.00135899054272
Gc3_35 0 n6 ns35 0 -0.00183705540269
Gc3_36 0 n6 ns36 0 0.00327369167124
Gc3_37 0 n6 ns37 0 -0.000823785381442
Gc3_38 0 n6 ns38 0 0.00248720657534
Gc3_39 0 n6 ns39 0 -0.000598023039958
Gc3_40 0 n6 ns40 0 -0.000107654172629
Gc3_41 0 n6 ns41 0 -0.00061898248816
Gc3_42 0 n6 ns42 0 0.000892397014269
Gc3_43 0 n6 ns43 0 0.000574020874682
Gc3_44 0 n6 ns44 0 -2.64430416307e-006
Gc3_45 0 n6 ns45 0 -0.0593383198323
Gc3_46 0 n6 ns46 0 -0.0735828516722
Gc3_47 0 n6 ns47 0 0.00622363336467
Gc3_48 0 n6 ns48 0 -0.0130071314472
Gc3_49 0 n6 ns49 0 -0.00995628444817
Gc3_50 0 n6 ns50 0 -0.00605491706667
Gc3_51 0 n6 ns51 0 -0.00102526907966
Gc3_52 0 n6 ns52 0 4.06599683626e-005
Gc3_53 0 n6 ns53 0 -8.87905359305e-005
Gc3_54 0 n6 ns54 0 2.06682954552e-005
Gc3_55 0 n6 ns55 0 -0.00317509459669
Gc3_56 0 n6 ns56 0 0.00323250156007
Gc3_57 0 n6 ns57 0 -0.00525374750053
Gc3_58 0 n6 ns58 0 -0.00147598862992
Gc3_59 0 n6 ns59 0 -0.00339118904103
Gc3_60 0 n6 ns60 0 0.00291773911587
Gc3_61 0 n6 ns61 0 -0.00115957912504
Gc3_62 0 n6 ns62 0 -0.0033090322364
Gc3_63 0 n6 ns63 0 -0.0010444280023
Gc3_64 0 n6 ns64 0 -0.00273127822918
Gc3_65 0 n6 ns65 0 -0.00107546381708
Gc3_66 0 n6 ns66 0 -0.00136240183917
Gc3_67 0 n6 ns67 0 0.0286948333406
Gc3_68 0 n6 ns68 0 0.0268324979238
Gc3_69 0 n6 ns69 0 0.00666047134928
Gc3_70 0 n6 ns70 0 0.0111231854313
Gc3_71 0 n6 ns71 0 -0.00268802713551
Gc3_72 0 n6 ns72 0 0.0031470075387
Gc3_73 0 n6 ns73 0 0.00128456529825
Gc3_74 0 n6 ns74 0 0.00203281356196
Gc3_75 0 n6 ns75 0 -4.59889921531e-005
Gc3_76 0 n6 ns76 0 6.25999851261e-006
Gc3_77 0 n6 ns77 0 -0.00275326905367
Gc3_78 0 n6 ns78 0 -0.00424377561213
Gc3_79 0 n6 ns79 0 0.00150842420655
Gc3_80 0 n6 ns80 0 -0.000663267836694
Gc3_81 0 n6 ns81 0 0.00251618399354
Gc3_82 0 n6 ns82 0 -0.00138435567206
Gc3_83 0 n6 ns83 0 0.00130824862215
Gc3_84 0 n6 ns84 0 0.0025095494155
Gc3_85 0 n6 ns85 0 0.0012845457475
Gc3_86 0 n6 ns86 0 0.000462926036445
Gc3_87 0 n6 ns87 0 -0.000705758174556
Gc3_88 0 n6 ns88 0 0.00152099822198
Gd3_1 0 n6 ni1 0 0.00415288714196
Gd3_2 0 n6 ni2 0 0.00561741499607
Gd3_3 0 n6 ni3 0 -0.0178815190119
Gd3_4 0 n6 ni4 0 0.00902490379672
Gc4_1 0 n8 ns1 0 0.0144285582063
Gc4_2 0 n8 ns2 0 0.00682394470379
Gc4_3 0 n8 ns3 0 0.00873922939655
Gc4_4 0 n8 ns4 0 0.00473349748016
Gc4_5 0 n8 ns5 0 0.000669887449411
Gc4_6 0 n8 ns6 0 -0.0002870801197
Gc4_7 0 n8 ns7 0 0.00207630136286
Gc4_8 0 n8 ns8 0 0.00280102908977
Gc4_9 0 n8 ns9 0 5.72424579871e-005
Gc4_10 0 n8 ns10 0 -1.01552806319e-005
Gc4_11 0 n8 ns11 0 0.00465884824921
Gc4_12 0 n8 ns12 0 0.00283977755579
Gc4_13 0 n8 ns13 0 -0.00162372104665
Gc4_14 0 n8 ns14 0 0.00026550482306
Gc4_15 0 n8 ns15 0 0.000596953459254
Gc4_16 0 n8 ns16 0 0.00283885421187
Gc4_17 0 n8 ns17 0 -0.000919828419142
Gc4_18 0 n8 ns18 0 4.78347385061e-005
Gc4_19 0 n8 ns19 0 -0.000878261185386
Gc4_20 0 n8 ns20 0 0.000758560274352
Gc4_21 0 n8 ns21 0 0.000637116922194
Gc4_22 0 n8 ns22 0 -0.000450429971812
Gc4_23 0 n8 ns23 0 -0.00780074486337
Gc4_24 0 n8 ns24 0 0.00696197514461
Gc4_25 0 n8 ns25 0 0.00571476170245
Gc4_26 0 n8 ns26 0 0.00685423150301
Gc4_27 0 n8 ns27 0 0.00935478104232
Gc4_28 0 n8 ns28 0 -0.00120210343955
Gc4_29 0 n8 ns29 0 -0.00215374306384
Gc4_30 0 n8 ns30 0 -0.0027767336754
Gc4_31 0 n8 ns31 0 5.95976813689e-005
Gc4_32 0 n8 ns32 0 -6.0584804425e-006
Gc4_33 0 n8 ns33 0 0.00182600250151
Gc4_34 0 n8 ns34 0 0.00246507442796
Gc4_35 0 n8 ns35 0 0.00442303691073
Gc4_36 0 n8 ns36 0 0.00346857391896
Gc4_37 0 n8 ns37 0 -0.000876197517794
Gc4_38 0 n8 ns38 0 0.00123412447969
Gc4_39 0 n8 ns39 0 -0.000302941381168
Gc4_40 0 n8 ns40 0 -0.00125495597139
Gc4_41 0 n8 ns41 0 -0.000955712963674
Gc4_42 0 n8 ns42 0 0.00241774336134
Gc4_43 0 n8 ns43 0 -0.000377749171731
Gc4_44 0 n8 ns44 0 0.0006457138437
Gc4_45 0 n8 ns45 0 0.0286976450791
Gc4_46 0 n8 ns46 0 0.0268259853463
Gc4_47 0 n8 ns47 0 0.00666906797481
Gc4_48 0 n8 ns48 0 0.0111247571811
Gc4_49 0 n8 ns49 0 -0.00268727380411
Gc4_50 0 n8 ns50 0 0.00315199090889
Gc4_51 0 n8 ns51 0 0.00129174333478
Gc4_52 0 n8 ns52 0 0.00203871573561
Gc4_53 0 n8 ns53 0 -4.6020247808e-005
Gc4_54 0 n8 ns54 0 6.41465603227e-006
Gc4_55 0 n8 ns55 0 -0.00277311464619
Gc4_56 0 n8 ns56 0 -0.00421280410236
Gc4_57 0 n8 ns57 0 0.00149744799758
Gc4_58 0 n8 ns58 0 -0.000672982094246
Gc4_59 0 n8 ns59 0 0.00250952235138
Gc4_60 0 n8 ns60 0 -0.00138652910401
Gc4_61 0 n8 ns61 0 0.00130991812408
Gc4_62 0 n8 ns62 0 0.002503872233
Gc4_63 0 n8 ns63 0 0.00128273049778
Gc4_64 0 n8 ns64 0 0.000454602409393
Gc4_65 0 n8 ns65 0 -0.000703784510173
Gc4_66 0 n8 ns66 0 0.0015222456204
Gc4_67 0 n8 ns67 0 -0.0364478084663
Gc4_68 0 n8 ns68 0 -0.0425185168063
Gc4_69 0 n8 ns69 0 0.00466461384306
Gc4_70 0 n8 ns70 0 -0.00478771843757
Gc4_71 0 n8 ns71 0 -0.0111793147288
Gc4_72 0 n8 ns72 0 -0.00296016517041
Gc4_73 0 n8 ns73 0 -0.00200233213205
Gc4_74 0 n8 ns74 0 -0.0014011060539
Gc4_75 0 n8 ns75 0 -7.9543820724e-005
Gc4_76 0 n8 ns76 0 1.47684765654e-005
Gc4_77 0 n8 ns77 0 -0.00019804760673
Gc4_78 0 n8 ns78 0 0.000306421255309
Gc4_79 0 n8 ns79 0 -0.00468232038902
Gc4_80 0 n8 ns80 0 0.000430738353135
Gc4_81 0 n8 ns81 0 -0.00113654214409
Gc4_82 0 n8 ns82 0 0.0021601158761
Gc4_83 0 n8 ns83 0 -0.000573907844554
Gc4_84 0 n8 ns84 0 -0.00151345063785
Gc4_85 0 n8 ns85 0 -0.00153726254936
Gc4_86 0 n8 ns86 0 -0.00193858814605
Gc4_87 0 n8 ns87 0 -0.000645229914007
Gc4_88 0 n8 ns88 0 -0.00031302218305
Gd4_1 0 n8 ni1 0 0.00472690430176
Gd4_2 0 n8 ni2 0 0.00338809736277
Gd4_3 0 n8 ni3 0 0.00901055490318
Gd4_4 0 n8 ni4 0 -0.0156575865921
.ends
*$
* BEGIN ANSOFT HEADER
* node 1    Port1
* node 2    Port2
* node 3    Port3
* node 4    Port4
*  Project: Project10
*   Format: PSpice
*   Topckt: s748030024_sp
*     Date: Fri Sep 11 16:42:50 2020
*    Notes: Frequency range: 1e+007 to 1e+010 Hz, 1000 points
*         : Maximum number of poles: 10000
*         : S-Matrix fitting error tolerance: 0.005
*         : Causality check tolerance: auto
*         : Passivity enforcement: off
*         : Causality enforcement: off
*         : Fitting method: TWA
*         : Matrix fitting: By entire matrix
*         : Ensure Z-parameter accuracy: on
*         : Relative error control: off
*         : Common ground option: on
*         : Final fitting error: 0.103285
*         : Final model order: 40
* END ANSOFT HEADER

.subckt WE-CCMF_748030024 1 4 2 3
Vam1 1 n2 dc 0
Rport1 n2 0 50
Vam2 2 n4 dc 0
Rport2 n4 0 50
Vam3 3 n6 dc 0
Rport3 n6 0 50
Vam4 4 n8 dc 0
Rport4 n8 0 50

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1
Fi3 0 ni3 Vam3 50
Gi3 0 ni3 3 0 1
Rt3 ni3 0 1
Fi4 0 ni4 Vam4 50
Gi4 0 ni4 4 0 1
Rt4 ni4 0 1

Ca1 ns1 0 1e-012
Ca2 ns2 0 1e-012
Ra1 ns1 0 196.057879393
Ra2 ns2 0 196.057879393
Ga1 ns1 0 ns2 0 -0.00906136858812
Ga2 ns2 0 ns1 0 0.00906136858812
Ca3 ns3 0 1e-012
Ca4 ns4 0 1e-012
Ra3 ns3 0 70.5014537058
Ra4 ns4 0 70.5014537058
Ga3 ns3 0 ns4 0 -0.0196146706844
Ga4 ns4 0 ns3 0 0.0196146706844
Ca5 ns5 0 1e-012
Ca6 ns6 0 1e-012
Ra5 ns5 0 79.3029027028
Ra6 ns6 0 79.3029027028
Ga5 ns5 0 ns6 0 -0.0395669021713
Ga6 ns6 0 ns5 0 0.0395669021713
Ca7 ns7 0 1e-012
Ca8 ns8 0 1e-012
Ra7 ns7 0 1026.61532806
Ra8 ns8 0 1026.61532806
Ga7 ns7 0 ns8 0 -0.0454193177237
Ga8 ns8 0 ns7 0 0.0454193177237
Ca9 ns9 0 1e-012
Ca10 ns10 0 1e-012
Ra9 ns9 0 92.1744418237
Ra10 ns10 0 92.1744418237
Ga9 ns9 0 ns10 0 -0.0571889056546
Ga10 ns10 0 ns9 0 0.0571889056546
Ca11 ns11 0 1e-012
Ca12 ns12 0 1e-012
Ra11 ns11 0 196.057879393
Ra12 ns12 0 196.057879393
Ga11 ns11 0 ns12 0 -0.00906136858812
Ga12 ns12 0 ns11 0 0.00906136858812
Ca13 ns13 0 1e-012
Ca14 ns14 0 1e-012
Ra13 ns13 0 70.5014537058
Ra14 ns14 0 70.5014537058
Ga13 ns13 0 ns14 0 -0.0196146706844
Ga14 ns14 0 ns13 0 0.0196146706844
Ca15 ns15 0 1e-012
Ca16 ns16 0 1e-012
Ra15 ns15 0 79.3029027028
Ra16 ns16 0 79.3029027028
Ga15 ns15 0 ns16 0 -0.0395669021713
Ga16 ns16 0 ns15 0 0.0395669021713
Ca17 ns17 0 1e-012
Ca18 ns18 0 1e-012
Ra17 ns17 0 1026.61532806
Ra18 ns18 0 1026.61532806
Ga17 ns17 0 ns18 0 -0.0454193177237
Ga18 ns18 0 ns17 0 0.0454193177237
Ca19 ns19 0 1e-012
Ca20 ns20 0 1e-012
Ra19 ns19 0 92.1744418237
Ra20 ns20 0 92.1744418237
Ga19 ns19 0 ns20 0 -0.0571889056546
Ga20 ns20 0 ns19 0 0.0571889056546
Ca21 ns21 0 1e-012
Ca22 ns22 0 1e-012
Ra21 ns21 0 196.057879393
Ra22 ns22 0 196.057879393
Ga21 ns21 0 ns22 0 -0.00906136858812
Ga22 ns22 0 ns21 0 0.00906136858812
Ca23 ns23 0 1e-012
Ca24 ns24 0 1e-012
Ra23 ns23 0 70.5014537058
Ra24 ns24 0 70.5014537058
Ga23 ns23 0 ns24 0 -0.0196146706844
Ga24 ns24 0 ns23 0 0.0196146706844
Ca25 ns25 0 1e-012
Ca26 ns26 0 1e-012
Ra25 ns25 0 79.3029027028
Ra26 ns26 0 79.3029027028
Ga25 ns25 0 ns26 0 -0.0395669021713
Ga26 ns26 0 ns25 0 0.0395669021713
Ca27 ns27 0 1e-012
Ca28 ns28 0 1e-012
Ra27 ns27 0 1026.61532806
Ra28 ns28 0 1026.61532806
Ga27 ns27 0 ns28 0 -0.0454193177237
Ga28 ns28 0 ns27 0 0.0454193177237
Ca29 ns29 0 1e-012
Ca30 ns30 0 1e-012
Ra29 ns29 0 92.1744418237
Ra30 ns30 0 92.1744418237
Ga29 ns29 0 ns30 0 -0.0571889056546
Ga30 ns30 0 ns29 0 0.0571889056546
Ca31 ns31 0 1e-012
Ca32 ns32 0 1e-012
Ra31 ns31 0 196.057879393
Ra32 ns32 0 196.057879393
Ga31 ns31 0 ns32 0 -0.00906136858812
Ga32 ns32 0 ns31 0 0.00906136858812
Ca33 ns33 0 1e-012
Ca34 ns34 0 1e-012
Ra33 ns33 0 70.5014537058
Ra34 ns34 0 70.5014537058
Ga33 ns33 0 ns34 0 -0.0196146706844
Ga34 ns34 0 ns33 0 0.0196146706844
Ca35 ns35 0 1e-012
Ca36 ns36 0 1e-012
Ra35 ns35 0 79.3029027028
Ra36 ns36 0 79.3029027028
Ga35 ns35 0 ns36 0 -0.0395669021713
Ga36 ns36 0 ns35 0 0.0395669021713
Ca37 ns37 0 1e-012
Ca38 ns38 0 1e-012
Ra37 ns37 0 1026.61532806
Ra38 ns38 0 1026.61532806
Ga37 ns37 0 ns38 0 -0.0454193177237
Ga38 ns38 0 ns37 0 0.0454193177237
Ca39 ns39 0 1e-012
Ca40 ns40 0 1e-012
Ra39 ns39 0 92.1744418237
Ra40 ns40 0 92.1744418237
Ga39 ns39 0 ns40 0 -0.0571889056546
Ga40 ns40 0 ns39 0 0.0571889056546

Gb1_1 ns1 0 ni1 0 0.0119323977363
Gb3_1 ns3 0 ni1 0 0.0298717292417
Gb5_1 ns5 0 ni1 0 0.0435856409986
Gb7_1 ns7 0 ni1 0 0.0454402079866
Gb9_1 ns9 0 ni1 0 0.0592470090122
Gb11_2 ns11 0 ni2 0 0.0119323977363
Gb13_2 ns13 0 ni2 0 0.0298717292417
Gb15_2 ns15 0 ni2 0 0.0435856409986
Gb17_2 ns17 0 ni2 0 0.0454402079866
Gb19_2 ns19 0 ni2 0 0.0592470090122
Gb21_3 ns21 0 ni3 0 0.0119323977363
Gb23_3 ns23 0 ni3 0 0.0298717292417
Gb25_3 ns25 0 ni3 0 0.0435856409986
Gb27_3 ns27 0 ni3 0 0.0454402079866
Gb29_3 ns29 0 ni3 0 0.0592470090122
Gb31_4 ns31 0 ni4 0 0.0119323977363
Gb33_4 ns33 0 ni4 0 0.0298717292417
Gb35_4 ns35 0 ni4 0 0.0435856409986
Gb37_4 ns37 0 ni4 0 0.0454402079866
Gb39_4 ns39 0 ni4 0 0.0592470090122

Gc1_1 0 n2 ns1 0 0.00827443729507
Gc1_2 0 n2 ns2 0 0.0105718336197
Gc1_3 0 n2 ns3 0 -0.0323946448638
Gc1_4 0 n2 ns4 0 -0.00718530743036
Gc1_5 0 n2 ns5 0 -0.00419651931046
Gc1_6 0 n2 ns6 0 -0.00822873441929
Gc1_7 0 n2 ns7 0 -0.000140439367629
Gc1_8 0 n2 ns8 0 -3.752946839e-005
Gc1_9 0 n2 ns9 0 -0.00196066161788
Gc1_10 0 n2 ns10 0 -0.00603064793702
Gc1_11 0 n2 ns11 0 0.0113325377752
Gc1_12 0 n2 ns12 0 0.00497408047365
Gc1_13 0 n2 ns13 0 0.0263499247867
Gc1_14 0 n2 ns14 0 0.0237011826153
Gc1_15 0 n2 ns15 0 -0.00737057980628
Gc1_16 0 n2 ns16 0 -0.000681869297365
Gc1_17 0 n2 ns17 0 8.57208996725e-005
Gc1_18 0 n2 ns18 0 -8.33302599927e-005
Gc1_19 0 n2 ns19 0 0.00122002123692
Gc1_20 0 n2 ns20 0 0.00837023740702
Gc1_21 0 n2 ns21 0 0.00723557696477
Gc1_22 0 n2 ns22 0 -0.00116630801645
Gc1_23 0 n2 ns23 0 0.00399502765434
Gc1_24 0 n2 ns24 0 -0.00612216175079
Gc1_25 0 n2 ns25 0 0.00933127770103
Gc1_26 0 n2 ns26 0 0.0082691455855
Gc1_27 0 n2 ns27 0 -0.000120144268182
Gc1_28 0 n2 ns28 0 -3.1122260051e-006
Gc1_29 0 n2 ns29 0 -0.00394634455854
Gc1_30 0 n2 ns30 0 0.00293682501457
Gc1_31 0 n2 ns31 0 0.00694367216828
Gc1_32 0 n2 ns32 0 0.00265569737877
Gc1_33 0 n2 ns33 0 -0.00804012167287
Gc1_34 0 n2 ns34 0 -0.00432511407254
Gc1_35 0 n2 ns35 0 -0.0053690041341
Gc1_36 0 n2 ns36 0 0.00415473345791
Gc1_37 0 n2 ns37 0 9.70814628266e-005
Gc1_38 0 n2 ns38 0 -7.62743134284e-005
Gc1_39 0 n2 ns39 0 0.000335618969677
Gc1_40 0 n2 ns40 0 -0.00486871534518
Gd1_1 0 n2 ni1 0 -0.0100802409167
Gd1_2 0 n2 ni2 0 0.00687313331598
Gd1_3 0 n2 ni3 0 0.00621711894339
Gd1_4 0 n2 ni4 0 -0.000595936200015
Gc2_1 0 n4 ns1 0 0.0113380109753
Gc2_2 0 n4 ns2 0 0.00497028772114
Gc2_3 0 n4 ns3 0 0.0263646454212
Gc2_4 0 n4 ns4 0 0.0237198781733
Gc2_5 0 n4 ns5 0 -0.00737065468879
Gc2_6 0 n4 ns6 0 -0.000675192036592
Gc2_7 0 n4 ns7 0 8.57545126957e-005
Gc2_8 0 n4 ns8 0 -8.3297773122e-005
Gc2_9 0 n4 ns9 0 0.00120858217865
Gc2_10 0 n4 ns10 0 0.00837115636756
Gc2_11 0 n4 ns11 0 0.00663207917813
Gc2_12 0 n4 ns12 0 0.0115899432883
Gc2_13 0 n4 ns13 0 -0.0306550872591
Gc2_14 0 n4 ns14 0 -0.00915755665949
Gc2_15 0 n4 ns15 0 -0.00210709468849
Gc2_16 0 n4 ns16 0 -0.0045579256312
Gc2_17 0 n4 ns17 0 -2.48851721971e-005
Gc2_18 0 n4 ns18 0 0.000116962968059
Gc2_19 0 n4 ns19 0 -0.00429170931073
Gc2_20 0 n4 ns20 0 -0.00475322685481
Gc2_21 0 n4 ns21 0 0.00691286773885
Gc2_22 0 n4 ns22 0 0.00188967359296
Gc2_23 0 n4 ns23 0 -0.00552396242701
Gc2_24 0 n4 ns24 0 -0.00433724262392
Gc2_25 0 n4 ns25 0 -0.00345316616088
Gc2_26 0 n4 ns26 0 0.00535839910392
Gc2_27 0 n4 ns27 0 4.29796611488e-005
Gc2_28 0 n4 ns28 0 -0.000156788745642
Gc2_29 0 n4 ns29 0 8.96814739919e-005
Gc2_30 0 n4 ns30 0 -0.003666101777
Gc2_31 0 n4 ns31 0 0.00661461259806
Gc2_32 0 n4 ns32 0 0.00339036658429
Gc2_33 0 n4 ns33 0 -0.0111894139647
Gc2_34 0 n4 ns34 0 -0.0091108117516
Gc2_35 0 n4 ns35 0 0.00667329160307
Gc2_36 0 n4 ns36 0 -0.00142363347024
Gc2_37 0 n4 ns37 0 -8.63065743492e-006
Gc2_38 0 n4 ns38 0 0.000142867677687
Gc2_39 0 n4 ns39 0 -0.00147155197554
Gc2_40 0 n4 ns40 0 0.000780425090323
Gd2_1 0 n4 ni1 0 0.0068698602196
Gd2_2 0 n4 ni2 0 -0.0137097166172
Gd2_3 0 n4 ni3 0 0.000366457096238
Gd2_4 0 n4 ni4 0 0.00413454492673
Gc3_1 0 n6 ns1 0 0.00723702363545
Gc3_2 0 n6 ns2 0 -0.00116651551077
Gc3_3 0 n6 ns3 0 0.00400472148349
Gc3_4 0 n6 ns4 0 -0.00612402588771
Gc3_5 0 n6 ns5 0 0.00932933456373
Gc3_6 0 n6 ns6 0 0.00827789796486
Gc3_7 0 n6 ns7 0 -0.000120168291872
Gc3_8 0 n6 ns8 0 -3.18385774536e-006
Gc3_9 0 n6 ns9 0 -0.00394905804139
Gc3_10 0 n6 ns10 0 0.00293291860988
Gc3_11 0 n6 ns11 0 0.00691309255951
Gc3_12 0 n6 ns12 0 0.00189008918035
Gc3_13 0 n6 ns13 0 -0.00552897932507
Gc3_14 0 n6 ns14 0 -0.00433367630973
Gc3_15 0 n6 ns15 0 -0.00345833091311
Gc3_16 0 n6 ns16 0 0.00535334789308
Gc3_17 0 n6 ns17 0 4.3058244992e-005
Gc3_18 0 n6 ns18 0 -0.000156736895102
Gc3_19 0 n6 ns19 0 9.06541482853e-005
Gc3_20 0 n6 ns20 0 -0.00366805524891
Gc3_21 0 n6 ns21 0 0.00925928276806
Gc3_22 0 n6 ns22 0 0.00798688152503
Gc3_23 0 n6 ns23 0 -0.0267660774488
Gc3_24 0 n6 ns24 0 -0.00626601080631
Gc3_25 0 n6 ns25 0 -0.000731535965374
Gc3_26 0 n6 ns26 0 -0.00755678039327
Gc3_27 0 n6 ns27 0 -7.14582692204e-005
Gc3_28 0 n6 ns28 0 9.77275536312e-005
Gc3_29 0 n6 ns29 0 -0.000962988130602
Gc3_30 0 n6 ns30 0 -0.00360234736809
Gc3_31 0 n6 ns31 0 0.010107847264
Gc3_32 0 n6 ns32 0 0.00604681261385
Gc3_33 0 n6 ns33 0 0.0233830055275
Gc3_34 0 n6 ns34 0 0.0204709428359
Gc3_35 0 n6 ns35 0 -0.00817101531568
Gc3_36 0 n6 ns36 0 -0.000380432515635
Gc3_37 0 n6 ns37 0 6.16184411032e-005
Gc3_38 0 n6 ns38 0 -9.21026281571e-005
Gc3_39 0 n6 ns39 0 0.00180685160109
Gc3_40 0 n6 ns40 0 0.00698324698169
Gd3_1 0 n6 ni1 0 0.00622002817608
Gd3_2 0 n6 ni2 0 0.000364039736222
Gd3_3 0 n6 ni3 0 -0.00514400997755
Gd3_4 0 n6 ni4 0 0.00588983758969
Gc4_1 0 n8 ns1 0 0.00694689627469
Gc4_2 0 n8 ns2 0 0.00265689347465
Gc4_3 0 n8 ns3 0 -0.00803344246832
Gc4_4 0 n8 ns4 0 -0.00432999632276
Gc4_5 0 n8 ns5 0 -0.00537272303639
Gc4_6 0 n8 ns6 0 0.00415273631928
Gc4_7 0 n8 ns7 0 9.71351160062e-005
Gc4_8 0 n8 ns8 0 -7.62116131592e-005
Gc4_9 0 n8 ns9 0 0.00034275029589
Gc4_10 0 n8 ns10 0 -0.00486784018089
Gc4_11 0 n8 ns11 0 0.00661931058903
Gc4_12 0 n8 ns12 0 0.00338708607407
Gc4_13 0 n8 ns13 0 -0.0111789850537
Gc4_14 0 n8 ns14 0 -0.00910992558827
Gc4_15 0 n8 ns15 0 0.0066775161667
Gc4_16 0 n8 ns16 0 -0.00141874190069
Gc4_17 0 n8 ns17 0 -8.81622854197e-006
Gc4_18 0 n8 ns18 0 0.000142906639511
Gc4_19 0 n8 ns19 0 -0.001471051705
Gc4_20 0 n8 ns20 0 0.000781571676441
Gc4_21 0 n8 ns21 0 0.0101013043623
Gc4_22 0 n8 ns22 0 0.00604916509816
Gc4_23 0 n8 ns23 0 0.0233762728652
Gc4_24 0 n8 ns24 0 0.0204745521727
Gc4_25 0 n8 ns25 0 -0.00818165570166
Gc4_26 0 n8 ns26 0 -0.000384183271732
Gc4_27 0 n8 ns27 0 6.15307217012e-005
Gc4_28 0 n8 ns28 0 -9.22461011585e-005
Gc4_29 0 n8 ns29 0 0.00180296760161
Gc4_30 0 n8 ns30 0 0.00697690485047
Gc4_31 0 n8 ns31 0 0.00903248244643
Gc4_32 0 n8 ns32 0 0.0102721086863
Gc4_33 0 n8 ns33 0 -0.0263918555748
Gc4_34 0 n8 ns34 0 -0.00862179791354
Gc4_35 0 n8 ns35 0 0.00175901038286
Gc4_36 0 n8 ns36 0 -0.00316796870082
Gc4_37 0 n8 ns37 0 -7.0714788761e-005
Gc4_38 0 n8 ns38 0 0.000143225005806
Gc4_39 0 n8 ns39 0 -0.00420755894251
Gc4_40 0 n8 ns40 0 -0.00222812858356
Gd4_1 0 n8 ni1 0 -0.000584932757019
Gd4_2 0 n8 ni2 0 0.00414273895197
Gd4_3 0 n8 ni3 0 0.00588036864334
Gd4_4 0 n8 ni4 0 -0.0100504535737
.ends
*$
* BEGIN ANSOFT HEADER
* node 1    Port1
* node 2    Port2
* node 3    Port3
* node 4    Port4
*  Project: Project10
*   Format: PSpice
*   Topckt: s748032455_sp
*     Date: Fri Sep 11 16:44:16 2020
*    Notes: Frequency range: 1e+007 to 1e+010 Hz, 1000 points
*         : Maximum number of poles: 10000
*         : S-Matrix fitting error tolerance: 0.005
*         : Causality check tolerance: auto
*         : Passivity enforcement: off
*         : Causality enforcement: off
*         : Fitting method: TWA
*         : Matrix fitting: By entire matrix
*         : Ensure Z-parameter accuracy: on
*         : Relative error control: off
*         : Common ground option: on
*         : Final fitting error: 0.147149
*         : Final model order: 32
* END ANSOFT HEADER

.subckt WE-CCMF_748032455 1 4 2 3
Vam1 1 n2 dc 0
Rport1 n2 0 50
Vam2 2 n4 dc 0
Rport2 n4 0 50
Vam3 3 n6 dc 0
Rport3 n6 0 50
Vam4 4 n8 dc 0
Rport4 n8 0 50

Fi1 0 ni1 Vam1 50
Gi1 0 ni1 1 0 1
Rt1 ni1 0 1
Fi2 0 ni2 Vam2 50
Gi2 0 ni2 2 0 1
Rt2 ni2 0 1
Fi3 0 ni3 Vam3 50
Gi3 0 ni3 3 0 1
Rt3 ni3 0 1
Fi4 0 ni4 Vam4 50
Gi4 0 ni4 4 0 1
Rt4 ni4 0 1

Ca1 ns1 0 1e-012
Ca2 ns2 0 1e-012
Ra1 ns1 0 137.905263418
Ra2 ns2 0 137.905263418
Ga1 ns1 0 ns2 0 -0.0114719812296
Ga2 ns2 0 ns1 0 0.0114719812296
Ca3 ns3 0 1e-012
Ca4 ns4 0 1e-012
Ra3 ns3 0 72.7955566495
Ra4 ns4 0 72.7955566495
Ga3 ns3 0 ns4 0 -0.0264867147809
Ga4 ns4 0 ns3 0 0.0264867147809
Ca5 ns5 0 1e-012
Ca6 ns6 0 1e-012
Ra5 ns5 0 131.988444403
Ra6 ns6 0 131.988444403
Ga5 ns5 0 ns6 0 -0.0412398646493
Ga6 ns6 0 ns5 0 0.0412398646493
Ca7 ns7 0 1e-012
Ca8 ns8 0 1e-012
Ra7 ns7 0 73.6333491313
Ra8 ns8 0 73.6333491313
Ga7 ns7 0 ns8 0 -0.057905345779
Ga8 ns8 0 ns7 0 0.057905345779
Ca9 ns9 0 1e-012
Ca10 ns10 0 1e-012
Ra9 ns9 0 137.905263418
Ra10 ns10 0 137.905263418
Ga9 ns9 0 ns10 0 -0.0114719812296
Ga10 ns10 0 ns9 0 0.0114719812296
Ca11 ns11 0 1e-012
Ca12 ns12 0 1e-012
Ra11 ns11 0 72.7955566495
Ra12 ns12 0 72.7955566495
Ga11 ns11 0 ns12 0 -0.0264867147809
Ga12 ns12 0 ns11 0 0.0264867147809
Ca13 ns13 0 1e-012
Ca14 ns14 0 1e-012
Ra13 ns13 0 131.988444403
Ra14 ns14 0 131.988444403
Ga13 ns13 0 ns14 0 -0.0412398646493
Ga14 ns14 0 ns13 0 0.0412398646493
Ca15 ns15 0 1e-012
Ca16 ns16 0 1e-012
Ra15 ns15 0 73.6333491313
Ra16 ns16 0 73.6333491313
Ga15 ns15 0 ns16 0 -0.057905345779
Ga16 ns16 0 ns15 0 0.057905345779
Ca17 ns17 0 1e-012
Ca18 ns18 0 1e-012
Ra17 ns17 0 137.905263418
Ra18 ns18 0 137.905263418
Ga17 ns17 0 ns18 0 -0.0114719812296
Ga18 ns18 0 ns17 0 0.0114719812296
Ca19 ns19 0 1e-012
Ca20 ns20 0 1e-012
Ra19 ns19 0 72.7955566495
Ra20 ns20 0 72.7955566495
Ga19 ns19 0 ns20 0 -0.0264867147809
Ga20 ns20 0 ns19 0 0.0264867147809
Ca21 ns21 0 1e-012
Ca22 ns22 0 1e-012
Ra21 ns21 0 131.988444403
Ra22 ns22 0 131.988444403
Ga21 ns21 0 ns22 0 -0.0412398646493
Ga22 ns22 0 ns21 0 0.0412398646493
Ca23 ns23 0 1e-012
Ca24 ns24 0 1e-012
Ra23 ns23 0 73.6333491313
Ra24 ns24 0 73.6333491313
Ga23 ns23 0 ns24 0 -0.057905345779
Ga24 ns24 0 ns23 0 0.057905345779
Ca25 ns25 0 1e-012
Ca26 ns26 0 1e-012
Ra25 ns25 0 137.905263418
Ra26 ns26 0 137.905263418
Ga25 ns25 0 ns26 0 -0.0114719812296
Ga26 ns26 0 ns25 0 0.0114719812296
Ca27 ns27 0 1e-012
Ca28 ns28 0 1e-012
Ra27 ns27 0 72.7955566495
Ra28 ns28 0 72.7955566495
Ga27 ns27 0 ns28 0 -0.0264867147809
Ga28 ns28 0 ns27 0 0.0264867147809
Ca29 ns29 0 1e-012
Ca30 ns30 0 1e-012
Ra29 ns29 0 131.988444403
Ra30 ns30 0 131.988444403
Ga29 ns29 0 ns30 0 -0.0412398646493
Ga30 ns30 0 ns29 0 0.0412398646493
Ca31 ns31 0 1e-012
Ca32 ns32 0 1e-012
Ra31 ns31 0 73.6333491313
Ra32 ns32 0 73.6333491313
Ga31 ns31 0 ns32 0 -0.057905345779
Ga32 ns32 0 ns31 0 0.057905345779

Gb1_1 ns1 0 ni1 0 0.0160555092211
Gb3_1 ns3 0 ni1 0 0.0336113422738
Gb5_1 ns5 0 ni1 0 0.042631773986
Gb7_1 ns7 0 ni1 0 0.0610905129583
Gb9_2 ns9 0 ni2 0 0.0160555092211
Gb11_2 ns11 0 ni2 0 0.0336113422738
Gb13_2 ns13 0 ni2 0 0.042631773986
Gb15_2 ns15 0 ni2 0 0.0610905129583
Gb17_3 ns17 0 ni3 0 0.0160555092211
Gb19_3 ns19 0 ni3 0 0.0336113422738
Gb21_3 ns21 0 ni3 0 0.042631773986
Gb23_3 ns23 0 ni3 0 0.0610905129583
Gb25_4 ns25 0 ni4 0 0.0160555092211
Gb27_4 ns27 0 ni4 0 0.0336113422738
Gb29_4 ns29 0 ni4 0 0.042631773986
Gb31_4 ns31 0 ni4 0 0.0610905129583

Gc1_1 0 n2 ns1 0 0.0163759606718
Gc1_2 0 n2 ns2 0 0.0060410177421
Gc1_3 0 n2 ns3 0 -0.0101830953862
Gc1_4 0 n2 ns4 0 -0.00303559015589
Gc1_5 0 n2 ns5 0 0.010060807327
Gc1_6 0 n2 ns6 0 0.0017993618469
Gc1_7 0 n2 ns7 0 -0.00542107660207
Gc1_8 0 n2 ns8 0 0.00468072312836
Gc1_9 0 n2 ns9 0 0.0165104213982
Gc1_10 0 n2 ns10 0 0.00654394319145
Gc1_11 0 n2 ns11 0 0.020655294427
Gc1_12 0 n2 ns12 0 0.018282647217
Gc1_13 0 n2 ns13 0 0.000744429962273
Gc1_14 0 n2 ns14 0 0.00263565251694
Gc1_15 0 n2 ns15 0 -0.00915557648611
Gc1_16 0 n2 ns16 0 0.00816361265957
Gc1_17 0 n2 ns17 0 0.0120001260226
Gc1_18 0 n2 ns18 0 -0.00334843428593
Gc1_19 0 n2 ns19 0 -0.00320017453016
Gc1_20 0 n2 ns20 0 2.74451083931e-005
Gc1_21 0 n2 ns21 0 0.00630611970698
Gc1_22 0 n2 ns22 0 -0.00168040769958
Gc1_23 0 n2 ns23 0 0.00363593878528
Gc1_24 0 n2 ns24 0 0.00425421977003
Gc1_25 0 n2 ns25 0 0.0109754352364
Gc1_26 0 n2 ns26 0 -0.00108363073468
Gc1_27 0 n2 ns27 0 -0.00386092026955
Gc1_28 0 n2 ns28 0 0.00169032348478
Gc1_29 0 n2 ns29 0 0.000752020574444
Gc1_30 0 n2 ns30 0 0.00162953486663
Gc1_31 0 n2 ns31 0 0.00122842609369
Gc1_32 0 n2 ns32 0 0.00294067903568
Gd1_1 0 n2 ni1 0 -0.00181674046838
Gd1_2 0 n2 ni2 0 0.00215954989418
Gd1_3 0 n2 ni3 0 0.0099080886979
Gd1_4 0 n2 ni4 0 0.00102517617064
Gc2_1 0 n4 ns1 0 0.0165125021765
Gc2_2 0 n4 ns2 0 0.00654680500644
Gc2_3 0 n4 ns3 0 0.0206549268088
Gc2_4 0 n4 ns4 0 0.0182861639603
Gc2_5 0 n4 ns5 0 0.000742612114314
Gc2_6 0 n4 ns6 0 0.0026353048325
Gc2_7 0 n4 ns7 0 -0.00915834554232
Gc2_8 0 n4 ns8 0 0.00816381131904
Gc2_9 0 n4 ns9 0 0.0101119872239
Gc2_10 0 n4 ns10 0 0.00938425794409
Gc2_11 0 n4 ns11 0 -0.0243404447362
Gc2_12 0 n4 ns12 0 0.0029808869958
Gc2_13 0 n4 ns13 0 0.00158800156115
Gc2_14 0 n4 ns14 0 -0.000367737162894
Gc2_15 0 n4 ns15 0 -0.00590687749443
Gc2_16 0 n4 ns16 0 -0.00415251659627
Gc2_17 0 n4 ns17 0 0.0113669879357
Gc2_18 0 n4 ns18 0 -0.00209134392696
Gc2_19 0 n4 ns19 0 -0.00115303184172
Gc2_20 0 n4 ns20 0 0.000805574050304
Gc2_21 0 n4 ns21 0 0.0021481817679
Gc2_22 0 n4 ns22 0 0.00214376550053
Gc2_23 0 n4 ns23 0 0.00168255672679
Gc2_24 0 n4 ns24 0 0.0047483340738
Gc2_25 0 n4 ns25 0 0.00748645292094
Gc2_26 0 n4 ns26 0 0.00223920691868
Gc2_27 0 n4 ns27 0 -0.0135430791358
Gc2_28 0 n4 ns28 0 0.0007503523917
Gc2_29 0 n4 ns29 0 0.0012937396973
Gc2_30 0 n4 ns30 0 0.000937412610374
Gc2_31 0 n4 ns31 0 -0.00184119557215
Gc2_32 0 n4 ns32 0 -0.00447466538019
Gd2_1 0 n4 ni1 0 0.00215590410319
Gd2_2 0 n4 ni2 0 -0.0233432722319
Gd2_3 0 n4 ni3 0 0.00269252278597
Gd2_4 0 n4 ni4 0 -0.00167966971907
Gc3_1 0 n6 ns1 0 0.0120068016928
Gc3_2 0 n6 ns2 0 -0.00335214629302
Gc3_3 0 n6 ns3 0 -0.00319713021974
Gc3_4 0 n6 ns4 0 3.21626451775e-005
Gc3_5 0 n6 ns5 0 0.00630673482663
Gc3_6 0 n6 ns6 0 -0.0016802991944
Gc3_7 0 n6 ns7 0 0.00363646912492
Gc3_8 0 n6 ns8 0 0.00425584043779
Gc3_9 0 n6 ns9 0 0.0113704185993
Gc3_10 0 n6 ns10 0 -0.00209270619742
Gc3_11 0 n6 ns11 0 -0.00115235931971
Gc3_12 0 n6 ns12 0 0.000809468915486
Gc3_13 0 n6 ns13 0 0.00214691269647
Gc3_14 0 n6 ns14 0 0.00214304838332
Gc3_15 0 n6 ns15 0 0.00168323686028
Gc3_16 0 n6 ns16 0 0.00474793363943
Gc3_17 0 n6 ns17 0 0.0158309230168
Gc3_18 0 n6 ns18 0 0.00669546985649
Gc3_19 0 n6 ns19 0 -0.0112057124689
Gc3_20 0 n6 ns20 0 -0.00417978159798
Gc3_21 0 n6 ns21 0 0.00963844848896
Gc3_22 0 n6 ns22 0 0.00182079491498
Gc3_23 0 n6 ns23 0 -0.00412581707681
Gc3_24 0 n6 ns24 0 0.00425528143529
Gc3_25 0 n6 ns25 0 0.0161038168044
Gc3_26 0 n6 ns26 0 0.00613425379329
Gc3_27 0 n6 ns27 0 0.021708011572
Gc3_28 0 n6 ns28 0 0.0166004200489
Gc3_29 0 n6 ns29 0 0.00250023382171
Gc3_30 0 n6 ns30 0 0.00333853225408
Gc3_31 0 n6 ns31 0 -0.00931626057888
Gc3_32 0 n6 ns32 0 0.00878717212091
Gd3_1 0 n6 ni1 0 0.00991185183934
Gd3_2 0 n6 ni2 0 0.00269373841587
Gd3_3 0 n6 ni3 0 -0.00134975577885
Gd3_4 0 n6 ni4 0 0.00372986450169
Gc4_1 0 n8 ns1 0 0.0109859425896
Gc4_2 0 n8 ns2 0 -0.0010870658907
Gc4_3 0 n8 ns3 0 -0.00385577661707
Gc4_4 0 n8 ns4 0 0.00169544555725
Gc4_5 0 n8 ns5 0 0.00075291278233
Gc4_6 0 n8 ns6 0 0.00163271360514
Gc4_7 0 n8 ns7 0 0.0012273294198
Gc4_8 0 n8 ns8 0 0.00294460471098
Gc4_9 0 n8 ns9 0 0.00749216340753
Gc4_10 0 n8 ns10 0 0.00223884186439
Gc4_11 0 n8 ns11 0 -0.0135457802023
Gc4_12 0 n8 ns12 0 0.000753185734976
Gc4_13 0 n8 ns13 0 0.001293637751
Gc4_14 0 n8 ns14 0 0.000937782237717
Gc4_15 0 n8 ns15 0 -0.00184114911193
Gc4_16 0 n8 ns16 0 -0.00447558975404
Gc4_17 0 n8 ns17 0 0.0161001523174
Gc4_18 0 n8 ns18 0 0.00613689777898
Gc4_19 0 n8 ns19 0 0.0217049795393
Gc4_20 0 n8 ns20 0 0.0166014288453
Gc4_21 0 n8 ns21 0 0.00249924911241
Gc4_22 0 n8 ns22 0 0.00333804874764
Gc4_23 0 n8 ns23 0 -0.00931956630649
Gc4_24 0 n8 ns24 0 0.00878440923794
Gc4_25 0 n8 ns25 0 0.00858837026407
Gc4_26 0 n8 ns26 0 0.0109210409471
Gc4_27 0 n8 ns27 0 -0.0268534493041
Gc4_28 0 n8 ns28 0 0.00149700570657
Gc4_29 0 n8 ns29 0 0.000765248523118
Gc4_30 0 n8 ns30 0 0.000249141088958
Gc4_31 0 n8 ns31 0 -0.00688126874059
Gc4_32 0 n8 ns32 0 -0.0049427298681
Gd4_1 0 n8 ni1 0 0.0010266231635
Gd4_2 0 n8 ni2 0 -0.00167862387423
Gd4_3 0 n8 ni3 0 0.00372546366711
Gd4_4 0 n8 ni4 0 -0.0256218701932
.ends
