**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 THT Power Inductor
* Matchcode:             WE-FAMI
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/9/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1012_744750340047_4.7u 1 2
Rp 1 2 2450
Cp 1 2 5.1p
Rs 1 N3 0.0066
L1 N3 2 4.5u
.ends 1012_744750340047_4.7u
*******
.subckt 1012_744750340150_15u 1 2
Rp 1 2 9250
Cp 1 2 9.6p
Rs 1 N3 0.0172
L1 N3 2 14u
.ends 1012_744750340150_15u
*******
.subckt 1215_744750460100_10u 1 2
Rp 1 2 3000
Cp 1 2 7.1p
Rs 1 N3 0.0067
L1 N3 2 9.5u
.ends 1215_744750460100_10u
*******
.subckt 1215_744750460150_15u 1 2
Rp 1 2 2160
Cp 1 2 22.3p
Rs 1 N3 0.0093
L1 N3 2 7u
.ends 1215_744750460150_15u
*******
.subckt 1215_744750460220_22u 1 2
Rp 1 2 5800
Cp 1 2 12.8p
Rs 1 N3 0.0124
L1 N3 2 18.5u
.ends 1215_744750460220_22u
*******
.subckt 1280_744750420047_4.7u 1 2
Rp 1 2 3120
Cp 1 2 7.2p
Rs 1 N3 0.007
L1 N3 2 5u
.ends 1280_744750420047_4.7u
*******
.subckt 1280_744750420068_6.8u 1 2
Rp 1 2 4000
Cp 1 2 6p
Rs 1 N3 0.0094
L1 N3 2 7u
.ends 1280_744750420068_6.8u
*******
.subckt 1280_744750420100_10u 1 2
Rp 1 2 5700
Cp 1 2 7.5p
Rs 1 N3 0.0129
L1 N3 2 10u
.ends 1280_744750420100_10u
*******
.subckt 1280_744750420150_15u 1 2
Rp 1 2 9500
Cp 1 2 6.6p
Rs 1 N3 0.0213
L1 N3 2 15u
.ends 1280_744750420150_15u
*******
.subckt 1280_744750420220_22u 1 2
Rp 1 2 13900
Cp 1 2 7.3p
Rs 1 N3 0.0309
L1 N3 2 23.5u
.ends 1280_744750420220_22u
*******
.subckt 1410_744750530047_4.7u 1 2
Rp 1 2 2500
Cp 1 2 9.35p
Rs 1 N3 0.0041
L1 N3 2 4.5u
.ends 1410_744750530047_4.7u
*******
.subckt 1410_744750530068_6.8u 1 2
Rp 1 2 3300
Cp 1 2 9.45p
Rs 1 N3 0.0053
L1 N3 2 6u
.ends 1410_744750530068_6.8u
*******
.subckt 1410_744750530100_10u 1 2
Rp 1 2 5450
Cp 1 2 11.1p
Rs 1 N3 0.008
L1 N3 2 10u
.ends 1410_744750530100_10u
*******
.subckt 1415_744750560047_4.7u 1 2
Rp 1 2 1300
Cp 1 2 5.95p
Rs 1 N3 0.0031
L1 N3 2 4u
.ends 1415_744750560047_4.7u
*******
.subckt 1415_744750560100_10u 1 2
Rp 1 2 3350
Cp 1 2 11.85p
Rs 1 N3 0.0054
L1 N3 2 10u
.ends 1415_744750560100_10u
*******
.subckt 1415_744750560220_22u 1 2
Rp 1 2 6800
Cp 1 2 14.25003492402p
Rs 1 N3 0.0126
L1 N3 2 23u
.ends 1415_744750560220_22u
*******
.subckt 8010_744750230030_3u 1 2
Rp 1 2 1560
Cp 1 2 2.94p
Rs 1 N3 0.007
L1 N3 2 3u
.ends 8010_744750230030_3u
*******
.subckt 8010_744750230047_4.7u 1 2
Rp 1 2 2720
Cp 1 2 4.4p
Rs 1 N3 0.0097
L1 N3 2 4.5u
.ends 8010_744750230047_4.7u
*******
.subckt 8010_744750230068_6.8u 1 2
Rp 1 2 3920
Cp 1 2 6.6p
Rs 1 N3 0.0122
L1 N3 2 6.5u
.ends 8010_744750230068_6.8u
*******
.subckt 8010_744750230100_10u 1 2
Rp 1 2 4900
Cp 1 2 7.7p
Rs 1 N3 0.0186
L1 N3 2 9.5u
.ends 8010_744750230100_10u
*******
.subckt 8010_744750230150_15u 1 2
Rp 1 2 7200
Cp 1 2 9.3p
Rs 1 N3 0.0279
L1 N3 2 14.5u
.ends 8010_744750230150_15u
*******
