**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  PFC Chokes
* Matchcode:              WE-PFC
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Toby      
* Date and Time:          2022-05-17
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt WE_PFC  1  2  3  4  PARAMS:
+  Lp=1
+  C=1
+  Rparp=1
+  Rserp=1
+  Cparp=1
+  Rsers=1
+  Ls=1
+  Cpars=1
+  Rpars=1
+  K=1
L_L1  1  N00180  {Lp}
C_C1  2  4  {C}  TC=0,0  
R_R50  2  4  1000g
C_C2  3  1  {C}  TC=0,0
R_R1  1  2  {Rparp}  TC=0,0
R_R2  N00180  2  {Rserp}  TC=0,0
C_C3  1  2  {Cparp}  TC=0,0
R_R3  N00984  4  {Rsers}  TC=0,0
L_L2  3  N00984  {Ls}
C_C4  3  4  {Cpars}  TC=0,0
R_R4  3  4  {Rpars}  TC=0,0
Kn_K1  L_L1  L_L2  {K}  
.ends  WE_PFC
  
.subckt 760800080  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00176681
+  C=.00000000001385
+  Rparp=2310
+  Rserp=1.3511
+  Cparp=.00000000003889
+  Rsers=1.0058
+  Ls=.00001055
+  Cpars=.00000000647
+  Rpars=1659.02
+  K=.967727
.ends  
  
.subckt 760801130  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.0007576
+  C=.00000000001602
+  Rparp=2140
+  Rserp=.5541
+  Cparp=.00000000003642
+  Rsers=.24489
+  Ls=.000617
+  Cpars=.00000000457
+  Rpars=4281
+  K=.960251
.ends  
  
.subckt 760801131  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.0007874
+  C=.00000000001933
+  Rparp=1940
+  Rserp=.72
+  Cparp=.00000000003218
+  Rsers=.4162
+  Ls=.0000063
+  Cpars=.00000000553
+  Rpars=1384
+  K=.964818
.ends  
  
.subckt 760801030  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00066458
+  C=.00000000001527
+  Rparp=2210
+  Rserp=.3821
+  Cparp=.00000000003558
+  Rsers=.216
+  Ls=.00000595
+  Cpars=.0000000042
+  Rpars=2965
+  K=.956311
.ends  
  
.subckt 760801031  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00068081
+  C=.00000000001702
+  Rparp=2050
+  Rserp=.8036
+  Cparp=.00000000002304
+  Rsers=.3255
+  Ls=.00000538
+  Cpars=.00000000425
+  Rpars=1645
+  K=.971223
.ends  
  
.subckt 760801020  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00050026
+  C=.00000000001222
+  Rparp=1990
+  Rserp=.3054
+  Cparp=.00000000003003
+  Rsers=.15405
+  Ls=.00000355
+  Cpars=.00000000441
+  Rpars=1872
+  K=.958927
.ends  
  
.subckt 760801021  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00050143
+  C=.00000000001824
+  Rparp=1980
+  Rserp=.4467
+  Cparp=.00000000005055
+  Rsers=.3827
+  Ls=.00000469
+  Cpars=.0000000000562
+  Rpars=1062
+  K=.954648
.ends  
  
.subckt 760802122  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00046626
+  C=.00000000001304
+  Rparp=2810
+  Rserp=.27809
+  Cparp=.0000000000613
+  Rsers=.17045
+  Ls=.00000454
+  Cpars=.0000000063
+  Rpars=2350
+  K=.97466
.ends  
  
.subckt 760802112  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00037744
+  C=.00000000001196
+  Rparp=2160
+  Rserp=.30401
+  Cparp=.00000000003823
+  Rsers=.1521
+  Ls=.00000262
+  Cpars=.00000000557
+  Rpars=1001
+  K=.949205
.ends  
  
.subckt 760802113  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00034101
+  C=.00000000001475
+  Rparp=2560
+  Rserp=.3389
+  Cparp=.00000000005251
+  Rsers=.27934
+  Ls=.00000321
+  Cpars=.00000000628
+  Rpars=739.9
+  K=.950691
.ends  
  
.subckt 760803200  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00014896
+  C=.00000000001678
+  Rparp=2010
+  Rserp=.09613
+  Cparp=.00000000005854
+  Rsers=.12527
+  Ls=.00000155
+  Cpars=.00000000577
+  Rpars=341.5
+  K=.911202
.ends  
  
.subckt 760804310  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00031283
+  C=.00000000001428
+  Rparp=3150
+  Rserp=.14554
+  Cparp=.00000000004103
+  Rsers=.20223
+  Ls=.00000289
+  Cpars=.00000000438
+  Rpars=853.1
+  K=.942485
.ends  
  
.subckt 760804110  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00024844
+  C=.00000000001316
+  Rparp=2320
+  Rserp=.12958
+  Cparp=.00000000003561
+  Rsers=.16091
+  Ls=.00000329
+  Cpars=.00000000289
+  Rpars=1222
+  K=.958547
.ends  
  
.subckt 760804111  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00025784
+  C=.00000000001314
+  Rparp=2260
+  Rserp=.2013
+  Cparp=.00000000005112
+  Rsers=.2331
+  Ls=.00000257
+  Cpars=.00000000535
+  Rpars=435.7
+  K=.943834
.ends  
  
.subckt 760805410  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00022969
+  C=.00000000000972
+  Rparp=2370
+  Rserp=.07171
+  Cparp=.00000000004843
+  Rsers=.17955
+  Ls=.00000246
+  Cpars=.00000000468
+  Rpars=478.2
+  K=.935882
.ends  
  
.subckt 760805210  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00019857
+  C=.0000000001441
+  Rparp=2300
+  Rserp=.10177
+  Cparp=.00000000004248
+  Rsers=.18134
+  Ls=.00000334
+  Cpars=.00000000267
+  Rpars=1028
+  K=.959102
.ends  
  
.subckt 760805211  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00019974
+  C=.0000000001386
+  Rparp=2040
+  Rserp=.20364
+  Cparp=.00000000005479
+  Rsers=.23377
+  Ls=.000002206
+  Cpars=.00000000548
+  Rpars=399.6
+  K=.930631
.ends  
  
.subckt 760806302  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00031264
+  C=.00000000000722
+  Rparp=2450
+  Rserp=.14904
+  Cparp=.00000000001391
+  Rsers=.24629
+  Ls=.0000045
+  Cpars=.0000000011
+  Rpars=1762
+  K=.932417
.ends  
  
.subckt 760806400  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00018315
+  C=.00000000000875
+  Rparp=2710
+  Rserp=.05775
+  Cparp=.00000000004635
+  Rsers=.15327
+  Ls=.00000229
+  Cpars=.00000000381
+  Rpars=442.8
+  K=.937116
.ends  
  
.subckt 760806200  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00015556
+  C=.0000000000067
+  Rparp=2430
+  Rserp=.06869
+  Cparp=.00000000003238
+  Rsers=.15755
+  Ls=.00000233
+  Cpars=.00000000223
+  Rpars=614.3
+  K=.941732
.ends  
  
.subckt 760806201  1  2  3  4
X1  1  2  3  4  WE_PFC  PARAMS:
+  Lp=.00015026
+  C=.0000000000118
+  Rparp=2440
+  Rserp=.12308
+  Cparp=.00000000005084
+  Rsers=.24326
+  Ls=.000224
+  Cpars=.00000000477
+  Rpars=440.7
+  K=.939009
.ends  
  
  
  
