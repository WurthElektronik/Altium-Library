**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Polymer Capacitors
* Matchcode:             WCAP-PTG5
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 870025174001_180uF 1 2
Rser 1 3 0.006905501311
Lser 2 4 4.094243353E-09
C1 3 4 0.00018
Rpar 3 4 27777.7777777778
.ends 870025174001_180uF
*******
.subckt 870025174002_220uF 1 2
Rser 1 3 0.0093716159468
Lser 2 4 9.602062072E-09
C1 3 4 0.00022
Rpar 3 4 22743.6823104693
.ends 870025174002_220uF
*******
.subckt 870025174003_270uF 1 2
Rser 1 3 0.0097
Lser 2 4 0.0000000075
C1 3 4 0.00027
Rpar 3 4 18518.5185185185
.ends 870025174003_270uF
*******
.subckt 870025174004_330uF 1 2
Rser 1 3 0.00716837313604
Lser 2 4 4.679096856E-09
C1 3 4 0.00033
Rpar 3 4 15144.2307692308
.ends 870025174004_330uF
*******
.subckt 870025174005_390uF 1 2
Rser 1 3 0.00797415030085
Lser 2 4 4.37816718E-09
C1 3 4 0.00039
Rpar 3 4 12830.9572301426
.ends 870025174005_390uF
*******
.subckt 870025174006_470uF 1 2
Rser 1 3 0.0111157582576
Lser 2 4 4.86795439E-09
C1 3 4 0.00047
Rpar 3 4 10641.8918918919
.ends 870025174006_470uF
*******
.subckt 870025174007_560uF 1 2
Rser 1 3 0.0075521170177
Lser 2 4 5.334109962E-09
C1 3 4 0.00056
Rpar 3 4 8928.57142857143
.ends 870025174007_560uF
*******
.subckt 870025174008_680uF 1 2
Rser 1 3 0.00819443523404
Lser 2 4 4.570175049E-09
C1 3 4 0.00068
Rpar 3 4 14719.6261682243
.ends 870025174008_680uF
*******
.subckt 870025174009_820uF 1 2
Rser 1 3 0.00806382896647
Lser 2 4 4.372780952E-09
C1 3 4 0.00082
Rpar 3 4 12195.1219512195
.ends 870025174009_820uF
*******
.subckt 870025174011_1.2mF 1 2
Rser 1 3 0.00721568441348
Lser 2 4 4.92965886E-09
C1 3 4 0.0012
Rpar 3 4 8333.33333333333
.ends 870025174011_1.2mF
*******
.subckt 870025175010_1mF 1 2
Rser 1 3 0.00924882437386
Lser 2 4 9.512821116E-09
C1 3 4 0.001
Rpar 3 4 10000
.ends 870025175010_1mF
*******
.subckt 870025175012_1.5mF 1 2
Rser 1 3 0.00634588646005
Lser 2 4 5.728059933E-09
C1 3 4 0.0015
Rpar 3 4 6666.66666666667
.ends 870025175012_1.5mF
*******
.subckt 870025175013_2mF 1 2
Rser 1 3 0.00742975126421
Lser 2 4 7.206422988E-09
C1 3 4 0.002
Rpar 3 4 5000
.ends 870025175013_2mF
*******
.subckt 870025374001_100uF 1 2
Rser 1 3 0.00745648767437
Lser 2 4 4.264724229E-09
C1 3 4 0.0001
Rpar 3 4 100000
.ends 870025374001_100uF
*******
.subckt 870025374002_180uF 1 2
Rser 1 3 0.0100625147214
Lser 2 4 3.253968873E-09
C1 3 4 0.00018
Rpar 3 4 55555.5555555556
.ends 870025374002_180uF
*******
.subckt 870025374003_220uF 1 2
Rser 1 3 0.00918402068331
Lser 2 4 4.136458108E-09
C1 3 4 0.00022
Rpar 3 4 45454.5454545455
.ends 870025374003_220uF
*******
.subckt 870025374004_270uF 1 2
Rser 1 3 0.00914436252619
Lser 2 4 5.21755114E-09
C1 3 4 0.00027
Rpar 3 4 37037.037037037
.ends 870025374004_270uF
*******
.subckt 870025374005_330uF 1 2
Rser 1 3 0.011754358369
Lser 2 4 6.654333686E-09
C1 3 4 0.00033
Rpar 3 4 30303.0303030303
.ends 870025374005_330uF
*******
.subckt 870025374006_390uF 1 2
Rser 1 3 0.00954956361983
Lser 2 4 7.308620963E-09
C1 3 4 0.00039
Rpar 3 4 25641.0256410256
.ends 870025374006_390uF
*******
.subckt 870025374007_470uF 1 2
Rser 1 3 0.00709347866327
Lser 2 4 3.81090008E-09
C1 3 4 0.00047
Rpar 3 4 21276.5957446809
.ends 870025374007_470uF
*******
.subckt 870025375008_560uF 1 2
Rser 1 3 0.00948072872021
Lser 2 4 7.310215468E-09
C1 3 4 0.00056
Rpar 3 4 17857.1428571429
.ends 870025375008_560uF
*******
.subckt 870025375009_680uF 1 2
Rser 1 3 0.00888268910394
Lser 2 4 6.307698388E-09
C1 3 4 0.00068
Rpar 3 4 16000
.ends 870025375009_680uF
*******
.subckt 870025375010_820uF 1 2
Rser 1 3 0.00986909381245
Lser 2 4 8.385939187E-09
C1 3 4 0.00082
Rpar 3 4 16000
.ends 870025375010_820uF
*******
.subckt 870025574001_39uF 1 2
Rser 1 3 0.0119171299228
Lser 2 4 5.715137189E-09
C1 3 4 0.000039
Rpar 3 4 128205.128205128
.ends 870025574001_39uF
*******
.subckt 870025574002_47uF 1 2
Rser 1 3 0.0145806474385
Lser 2 4 4.121035102E-09
C1 3 4 0.000047
Rpar 3 4 106382.978723404
.ends 870025574002_47uF
*******
.subckt 870025574003_68uF 1 2
Rser 1 3 0.0120548630548
Lser 2 4 3.165824999E-09
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 870025574003_68uF
*******
.subckt 870025574004_82uF 1 2
Rser 1 3 0.010634120178
Lser 2 4 3.870316506E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 870025574004_82uF
*******
.subckt 870025574005_100uF 1 2
Rser 1 3 0.0139699926404
Lser 2 4 4.541094258E-09
C1 3 4 0.0001
Rpar 3 4 50000
.ends 870025574005_100uF
*******
.subckt 870025575006_180uF 1 2
Rser 1 3 0.00906261574775
Lser 2 4 6.046315918E-09
C1 3 4 0.00018
Rpar 3 4 27777.7777777778
.ends 870025575006_180uF
*******
.subckt 870025575007_220uF 1 2
Rser 1 3 0.0106752654807
Lser 2 4 6.530197714E-09
C1 3 4 0.00022
Rpar 3 4 22727.2727272727
.ends 870025575007_220uF
*******
.subckt 870025575008_270uF 1 2
Rser 1 3 0.0076197123697
Lser 2 4 5.27318462E-09
C1 3 4 0.00027
Rpar 3 4 18518.5185185185
.ends 870025575008_270uF
*******
.subckt 870025575009_330uF 1 2
Rser 1 3 0.00918245851494
Lser 2 4 5.937013811E-09
C1 3 4 0.00033
Rpar 3 4 15151.5151515152
.ends 870025575009_330uF
*******
