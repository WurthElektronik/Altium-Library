**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Bi-color TOP LED Waterclear
* Matchcode:              WL-SMTW
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-15
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 3528_150141RB73100 1 2 3 4
D1 1 3 Red
.MODEL Red D
+ IS=411.95E-18
+ N=2.2440
+ RS=.34593
+ IKF=704.53E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 2 4 Blue
.MODEL Blue D
+ IS=18.482E-6
+ N=4.1460
+ RS=1.2885
+ IKF=1.1173E-12
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141RV73100 1 2 3 4
D1 1 3 Red
.MODEL Red D
+ IS=83.143E-15
+ N=2.7379
+ RS=.505
+ IKF=800.56E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 2 4 Green
.MODEL Green D
+ IS=10.000E-21
+ N=1.7773
+ RS=1.0008E-6
+ IKF=1.0196E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141YB73100 1 2 3 4
D1 1 3 Yellow
.MODEL Yellow D
+ IS=11.252E-18
+ N=2.1040
+ RS=.29401
+ IKF=654.99E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 2 4 Blue
.MODEL Blue D
+ IS=3.7408E-9
+ N=4.3687
+ RS=1.4814
+ IKF=43.812E-9
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141YV73100 1 2 3 4
D1 1 3 Yellow
.MODEL Yellow D
+ IS=83.143E-15
+ N=2.7379
+ RS=.505
+ IKF=800.56E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 2 4 BGreen
.MODEL BGreen D
+ IS=10.000E-21
+ N=1.7773
+ RS=1.0000E-6
+ IKF=1.0200E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141RY73110 1 2 3 4
D1 1 3 Red
.MODEL Red D
+ IS=27.459E-15
+ N=2.5610
+ RS=.45359
+ IKF=780.07E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 4 2 Yellow
.MODEL Yellow D
+ IS=10.000E-21
+ N=1.7773
+ RS=1.0000E-6
+ IKF=1.0200E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141SV73110 1 2 3 4
D1 1 3 SRed
.MODEL SRed D
+ IS=15.170E-15
+ N=2.4744
+ RS=.42996
+ IKF=764.57E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 4 2 BGreen
.MODEL BGreen D
+ IS=10.000E-21
+ N=1.7773
+ RS=1.0000E-6
+ IKF=1.0200E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********
.subckt 3528_150141YV73110 1 2 3 4
D1 1 3 Yellow
.MODEL Yellow D
+ IS=83.143E-15
+ N=2.7379
+ RS=.505
+ IKF=800.56E-6
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
D2 4 2 BGreen
.MODEL BGreen D
+ IS=10.000E-21
+ N=1.7773
+ RS=1.0000E-6
+ IKF=1.0200E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
**********

















































