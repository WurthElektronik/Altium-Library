**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Electrolytic Capacitors
* Matchcode:             WCAP-ATLI
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 860080272001_68uF 1 2
Rser 1 3 0.27
Lser 2 4 0.0000000008
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860080272001_68uF
*******
.subckt 860080272002_82uF 1 2
Rser 1 3 0.258
Lser 2 4 0.000000001
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860080272002_82uF
*******
.subckt 860080272003_100uF 1 2
Rser 1 3 0.275089565456
Lser 2 4 5.153371331E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860080272003_100uF
*******
.subckt 860080272004_120uF 1 2
Rser 1 3 0.23422092106
Lser 2 4 5.055647368E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860080272004_120uF
*******
.subckt 860080273005_150uF 1 2
Rser 1 3 0.13
Lser 2 4 0.0000000022
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860080273005_150uF
*******
.subckt 860080273006_180uF 1 2
Rser 1 3 0.112
Lser 2 4 0.000000003
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860080273006_180uF
*******
.subckt 860080273007_220uF 1 2
Rser 1 3 0.11
Lser 2 4 0.000000003
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860080273007_220uF
*******
.subckt 860080273008_270uF 1 2
Rser 1 3 0.073
Lser 2 4 0.000000005
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860080273008_270uF
*******
.subckt 860080274009_330uF 1 2
Rser 1 3 0.078
Lser 2 4 0.000000005
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080274009_330uF
*******
.subckt 860080274010_390uF 1 2
Rser 1 3 0.089398341136
Lser 2 4 6.224049891E-09
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860080274010_390uF
*******
.subckt 860080274011_470uF 1 2
Rser 1 3 0.062
Lser 2 4 0.000000004
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860080274011_470uF
*******
.subckt 860080274012_560uF 1 2
Rser 1 3 0.052
Lser 2 4 0.000000005
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860080274012_560uF
*******
.subckt 860080274013_680uF 1 2
Rser 1 3 0.0414120202352
Lser 2 4 5.46208746E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860080274013_680uF
*******
.subckt 860080274014_820uF 1 2
Rser 1 3 0.04955
Lser 2 4 9.701418903E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860080274014_820uF
*******
.subckt 860080274015_1mF 1 2
Rser 1 3 0.0326404317137
Lser 2 4 5.672271496E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860080274015_1mF
*******
.subckt 860080275016_1mF 1 2
Rser 1 3 0.029949417198
Lser 2 4 7.449639234E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860080275016_1mF
*******
.subckt 860080275017_1.2mF 1 2
Rser 1 3 0.0230954455149
Lser 2 4 7.276968742E-09
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860080275017_1.2mF
*******
.subckt 860080275018_1.5mF 1 2
Rser 1 3 0.0226721623818
Lser 2 4 6.758324858E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860080275018_1.5mF
*******
.subckt 860080275019_1.8mF 1 2
Rser 1 3 0.019576368231
Lser 2 4 5.729423625E-09
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860080275019_1.8mF
*******
.subckt 860080278020_2.2mF 1 2
Rser 1 3 0.0205
Lser 2 4 0.000000004
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860080278020_2.2mF
*******
.subckt 860080278021_2.7mF 1 2
Rser 1 3 0.0188167552074
Lser 2 4 6.649611745E-09
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860080278021_2.7mF
*******
.subckt 860080278022_3.3mF 1 2
Rser 1 3 0.0172782827262
Lser 2 4 9.274805991E-09
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860080278022_3.3mF
*******
.subckt 860080278023_3.9mF 1 2
Rser 1 3 0.014900169292
Lser 2 4 7.984603749E-09
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860080278023_3.9mF
*******
.subckt 860080278024_4.7mF 1 2
Rser 1 3 0.0118492505591
Lser 2 4 1.042591744E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860080278024_4.7mF
*******
.subckt 860080280025_5.6mF 1 2
Rser 1 3 0.0141833798798
Lser 2 4 1.6437430262E-08
C1 3 4 0.0056
Rpar 3 4 17857.1428571429
.ends 860080280025_5.6mF
*******
.subckt 860080280026_6.8mF 1 2
Rser 1 3 0.0174251442304
Lser 2 4 1.9094745655E-08
C1 3 4 0.0068
Rpar 3 4 14705.8823529412
.ends 860080280026_6.8mF
*******
.subckt 860080372001_47uF 1 2
Rser 1 3 0.297840944306
Lser 2 4 4.941640767E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860080372001_47uF
*******
.subckt 860080372002_56uF 1 2
Rser 1 3 0.195
Lser 2 4 0.000000002
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860080372002_56uF
*******
.subckt 860080372003_68uF 1 2
Rser 1 3 0.178
Lser 2 4 0.000000002
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860080372003_68uF
*******
.subckt 860080372004_82uF 1 2
Rser 1 3 0.155
Lser 2 4 0.000000002
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860080372004_82uF
*******
.subckt 860080373005_100uF 1 2
Rser 1 3 0.157
Lser 2 4 0.000000003
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860080373005_100uF
*******
.subckt 860080373006_120uF 1 2
Rser 1 3 0.095
Lser 2 4 0.000000005
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860080373006_120uF
*******
.subckt 860080373007_150uF 1 2
Rser 1 3 0.124
Lser 2 4 8.957276225E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860080373007_150uF
*******
.subckt 860080374008_180uF 1 2
Rser 1 3 0.07
Lser 2 4 0.000000007
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860080374008_180uF
*******
.subckt 860080374009_220uF 1 2
Rser 1 3 0.087
Lser 2 4 0.000000003
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860080374009_220uF
*******
.subckt 860080374010_270uF 1 2
Rser 1 3 0.080558187659
Lser 2 4 6.529043091E-09
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860080374010_270uF
*******
.subckt 860080374011_330uF 1 2
Rser 1 3 0.06
Lser 2 4 0.000000006
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080374011_330uF
*******
.subckt 860080374012_390uF 1 2
Rser 1 3 0.05
Lser 2 4 0.000000008
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860080374012_390uF
*******
.subckt 860080374013_470uF 1 2
Rser 1 3 0.05
Lser 2 4 0.000000006
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860080374013_470uF
*******
.subckt 860080374015_560uF 1 2
Rser 1 3 0.0308471653784
Lser 2 4 5.229199481E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860080374015_560uF
*******
.subckt 860080374016_680uF 1 2
Rser 1 3 0.0326214765496
Lser 2 4 6.573791844E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860080374016_680uF
*******
.subckt 860080375014_470uF 1 2
Rser 1 3 0.0415523159563
Lser 2 4 5.41345812E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860080375014_470uF
*******
.subckt 860080375017_680uF 1 2
Rser 1 3 0.0294526329507
Lser 2 4 5.280787034E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860080375017_680uF
*******
.subckt 860080375018_820uF 1 2
Rser 1 3 0.0260966112518
Lser 2 4 6.030426301E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860080375018_820uF
*******
.subckt 860080375019_1mF 1 2
Rser 1 3 0.0217042631628
Lser 2 4 6.405811171E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860080375019_1mF
*******
.subckt 860080375020_1.2mF 1 2
Rser 1 3 0.0240810352057
Lser 2 4 5.678491644E-09
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860080375020_1.2mF
*******
.subckt 860080375021_1.5mF 1 2
Rser 1 3 0.0173451240768
Lser 2 4 8.419259316E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860080375021_1.5mF
*******
.subckt 860080378022_1.5mF 1 2
Rser 1 3 0.0209812031156
Lser 2 4 8.562278737E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860080378022_1.5mF
*******
.subckt 860080378023_1.8mF 1 2
Rser 1 3 0.0202388612411
Lser 2 4 7.368635803E-09
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860080378023_1.8mF
*******
.subckt 860080378024_2.2mF 1 2
Rser 1 3 0.023
Lser 2 4 0.000000011
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860080378024_2.2mF
*******
.subckt 860080378025_2.7mF 1 2
Rser 1 3 0.0165541180762
Lser 2 4 8.7503083E-09
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860080378025_2.7mF
*******
.subckt 860080378026_3.3mF 1 2
Rser 1 3 0.0124077453606
Lser 2 4 1.0816855727E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860080378026_3.3mF
*******
.subckt 860080380027_3.9mF 1 2
Rser 1 3 0.0175032711726
Lser 2 4 1.6038532234E-08
C1 3 4 0.0039
Rpar 3 4 25641.0256410256
.ends 860080380027_3.9mF
*******
.subckt 860080380028_4.7mF 1 2
Rser 1 3 0.014352702648
Lser 2 4 1.5779304244E-08
C1 3 4 0.0047
Rpar 3 4 21276.5957446809
.ends 860080380028_4.7mF
*******
.subckt 860080472001_39uF 1 2
Rser 1 3 0.235
Lser 2 4 0.0000000017
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860080472001_39uF
*******
.subckt 860080472002_47uF 1 2
Rser 1 3 0.218
Lser 2 4 0.0000000015
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860080472002_47uF
*******
.subckt 860080472003_56uF 1 2
Rser 1 3 0.162
Lser 2 4 0.000000002
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860080472003_56uF
*******
.subckt 860080473004_68uF 1 2
Rser 1 3 0.155
Lser 2 4 0.0000000032
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860080473004_68uF
*******
.subckt 860080473005_82uF 1 2
Rser 1 3 0.115
Lser 2 4 0.000000004
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860080473005_82uF
*******
.subckt 860080473006_100uF 1 2
Rser 1 3 0.112
Lser 2 4 0.0000000181
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860080473006_100uF
*******
.subckt 860080473007_120uF 1 2
Rser 1 3 0.1
Lser 2 4 0.000000005
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860080473007_120uF
*******
.subckt 860080474008_150uF 1 2
Rser 1 3 0.067
Lser 2 4 0.000000009
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860080474008_150uF
*******
.subckt 860080474009_180uF 1 2
Rser 1 3 0.0664134347643
Lser 2 4 3.953854409E-09
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860080474009_180uF
*******
.subckt 860080474010_220uF 1 2
Rser 1 3 0.065
Lser 2 4 0.0000000065
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860080474010_220uF
*******
.subckt 860080474011_270uF 1 2
Rser 1 3 0.05
Lser 2 4 0.000000009
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860080474011_270uF
*******
.subckt 860080474012_330uF 1 2
Rser 1 3 0.047373566599
Lser 2 4 6.401102138E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080474012_330uF
*******
.subckt 860080474015_470uF 1 2
Rser 1 3 0.033
Lser 2 4 0.000000007
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860080474015_470uF
*******
.subckt 860080475013_330uF 1 2
Rser 1 3 0.0432003779907
Lser 2 4 5.24470864E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080475013_330uF
*******
.subckt 860080475014_390uF 1 2
Rser 1 3 0.0400219042267
Lser 2 4 6.780485429E-09
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860080475014_390uF
*******
.subckt 860080475016_470uF 1 2
Rser 1 3 0.0319983465212
Lser 2 4 7.329806924E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860080475016_470uF
*******
.subckt 860080475017_560uF 1 2
Rser 1 3 0.0258470596199
Lser 2 4 8.898873769E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860080475017_560uF
*******
.subckt 860080475018_680uF 1 2
Rser 1 3 0.0219731549032
Lser 2 4 7.356909243E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860080475018_680uF
*******
.subckt 860080475019_820uF 1 2
Rser 1 3 0.0185549226115
Lser 2 4 7.521817968E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860080475019_820uF
*******
.subckt 860080478020_1mF 1 2
Rser 1 3 0.0375210685203
Lser 2 4 7.247446143E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860080478020_1mF
*******
.subckt 860080478021_1.2mF 1 2
Rser 1 3 0.022096584594
Lser 2 4 5.778062454E-09
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860080478021_1.2mF
*******
.subckt 860080478022_1.5mF 1 2
Rser 1 3 0.0168950222213
Lser 2 4 7.715165619E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860080478022_1.5mF
*******
.subckt 860080478023_1.8mF 1 2
Rser 1 3 0.0145878986049
Lser 2 4 8.235918493E-09
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860080478023_1.8mF
*******
.subckt 860080478024_2.2mF 1 2
Rser 1 3 0.019
Lser 2 4 0.00000001
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860080478024_2.2mF
*******
.subckt 860080480025_2.7mF 1 2
Rser 1 3 0.0218263165021
Lser 2 4 1.7708955251E-08
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860080480025_2.7mF
*******
.subckt 860080480026_3.3mF 1 2
Rser 1 3 0.0150467943442
Lser 2 4 1.4018478991E-08
C1 3 4 0.0033
Rpar 3 4 30303.0303030303
.ends 860080480026_3.3mF
*******
.subckt 860080572001_33uF 1 2
Rser 1 3 0.18
Lser 2 4 0.0000000028
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860080572001_33uF
*******
.subckt 860080573002_39uF 1 2
Rser 1 3 0.178
Lser 2 4 0.000000004
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860080573002_39uF
*******
.subckt 860080573003_47uF 1 2
Rser 1 3 0.133
Lser 2 4 0.0000000074
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860080573003_47uF
*******
.subckt 860080573004_56uF 1 2
Rser 1 3 0.12
Lser 2 4 0.0000000055
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860080573004_56uF
*******
.subckt 860080573005_68uF 1 2
Rser 1 3 0.1
Lser 2 4 0.000000006
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860080573005_68uF
*******
.subckt 860080574006_82uF 1 2
Rser 1 3 0.078
Lser 2 4 0.0000000075
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860080574006_82uF
*******
.subckt 860080574007_100uF 1 2
Rser 1 3 0.11
Lser 2 4 0.0000000065
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860080574007_100uF
*******
.subckt 860080574008_120uF 1 2
Rser 1 3 0.078
Lser 2 4 0.000000008
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860080574008_120uF
*******
.subckt 860080574009_150uF 1 2
Rser 1 3 0.058
Lser 2 4 0.000000008
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860080574009_150uF
*******
.subckt 860080574010_180uF 1 2
Rser 1 3 0.055
Lser 2 4 0.000000008
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860080574010_180uF
*******
.subckt 860080574011_220uF 1 2
Rser 1 3 0.047
Lser 2 4 0.000000006
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860080574011_220uF
*******
.subckt 860080574014_330uF 1 2
Rser 1 3 0.0287590173672
Lser 2 4 6.792920841E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080574014_330uF
*******
.subckt 860080575012_220uF 1 2
Rser 1 3 0.0442034368615
Lser 2 4 7.087476406E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860080575012_220uF
*******
.subckt 860080575013_270uF 1 2
Rser 1 3 0.0349063605163
Lser 2 4 4.993830281E-09
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860080575013_270uF
*******
.subckt 860080575015_330uF 1 2
Rser 1 3 0.0270805237152
Lser 2 4 6.177668085E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080575015_330uF
*******
.subckt 860080575016_390uF 1 2
Rser 1 3 0.0286771540686
Lser 2 4 7.88677152E-09
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860080575016_390uF
*******
.subckt 860080575017_470uF 1 2
Rser 1 3 0.031
Lser 2 4 0.000000008
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860080575017_470uF
*******
.subckt 860080575018_560uF 1 2
Rser 1 3 0.0170249712893
Lser 2 4 6.42235943E-09
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860080575018_560uF
*******
.subckt 860080578019_680uF 1 2
Rser 1 3 0.0221147982109
Lser 2 4 6.80477786E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860080578019_680uF
*******
.subckt 860080578020_820uF 1 2
Rser 1 3 0.0175276884178
Lser 2 4 8.765114263E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860080578020_820uF
*******
.subckt 860080578021_1mF 1 2
Rser 1 3 0.017264868876
Lser 2 4 7.21169756E-09
C1 3 4 0.001
Rpar 3 4 100000
.ends 860080578021_1mF
*******
.subckt 860080578022_1.2mF 1 2
Rser 1 3 0.02028
Lser 2 4 1.4912959568E-08
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860080578022_1.2mF
*******
.subckt 860080578024_1.5mF 1 2
Rser 1 3 0.0120221062137
Lser 2 4 9.316172841E-09
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860080578024_1.5mF
*******
.subckt 860080580023_1.2mF 1 2
Rser 1 3 0.0167625300837
Lser 2 4 1.7515264075E-08
C1 3 4 0.0012
Rpar 3 4 83333.3333333333
.ends 860080580023_1.2mF
*******
.subckt 860080580025_1.5mF 1 2
Rser 1 3 0.0138822735555
Lser 2 4 1.5516670418E-08
C1 3 4 0.0015
Rpar 3 4 66666.6666666667
.ends 860080580025_1.5mF
*******
.subckt 860080580026_1.8mF 1 2
Rser 1 3 0.0160751430576
Lser 2 4 1.8110019627E-08
C1 3 4 0.0018
Rpar 3 4 55555.5555555556
.ends 860080580026_1.8mF
*******
.subckt 860080580027_2.2mF 1 2
Rser 1 3 0.0114207043994
Lser 2 4 1.4322505729E-08
C1 3 4 0.0022
Rpar 3 4 45454.5454545455
.ends 860080580027_2.2mF
*******
.subckt 860080581028_2.7mF 1 2
Rser 1 3 0.0164649533682
Lser 2 4 1.6504712212E-08
C1 3 4 0.0027
Rpar 3 4 37037.037037037
.ends 860080581028_2.7mF
*******
.subckt 860080672001_22uF 1 2
Rser 1 3 0.21
Lser 2 4 0.0000000053
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860080672001_22uF
*******
.subckt 860080673002_27uF 1 2
Rser 1 3 0.134
Lser 2 4 0.0000000055
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 860080673002_27uF
*******
.subckt 860080673003_33uF 1 2
Rser 1 3 0.316099278456
Lser 2 4 5.183810129E-09
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860080673003_33uF
*******
.subckt 860080673004_39uF 1 2
Rser 1 3 0.245
Lser 2 4 0.0000000023
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860080673004_39uF
*******
.subckt 860080674005_47uF 1 2
Rser 1 3 0.11
Lser 2 4 0.000000007
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860080674005_47uF
*******
.subckt 860080674006_56uF 1 2
Rser 1 3 0.084
Lser 2 4 0.000000009
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860080674006_56uF
*******
.subckt 860080674007_68uF 1 2
Rser 1 3 0.071
Lser 2 4 0.00000001
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860080674007_68uF
*******
.subckt 860080674008_82uF 1 2
Rser 1 3 0.072
Lser 2 4 0.00000001
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860080674008_82uF
*******
.subckt 860080674009_100uF 1 2
Rser 1 3 0.095
Lser 2 4 0.0000000192
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860080674009_100uF
*******
.subckt 860080674010_120uF 1 2
Rser 1 3 0.06
Lser 2 4 0.00000001
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860080674010_120uF
*******
.subckt 860080674013_180uF 1 2
Rser 1 3 0.0355511452069
Lser 2 4 6.091403394E-09
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860080674013_180uF
*******
.subckt 860080675011_120uF 1 2
Rser 1 3 0.0484646880905
Lser 2 4 6.551735953E-09
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860080675011_120uF
*******
.subckt 860080675012_150uF 1 2
Rser 1 3 0.0421844483567
Lser 2 4 6.059123487E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860080675012_150uF
*******
.subckt 860080675014_180uF 1 2
Rser 1 3 0.0328489863998
Lser 2 4 6.766316192E-09
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860080675014_180uF
*******
.subckt 860080675015_220uF 1 2
Rser 1 3 0.0336226338474
Lser 2 4 4.721797344E-09
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860080675015_220uF
*******
.subckt 860080675016_270uF 1 2
Rser 1 3 0.0263754087233
Lser 2 4 7.034767306E-09
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860080675016_270uF
*******
.subckt 860080675017_330uF 1 2
Rser 1 3 0.0238746414646
Lser 2 4 5.007853336E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080675017_330uF
*******
.subckt 860080678018_390uF 1 2
Rser 1 3 0.0235710491505
Lser 2 4 9.349354916E-09
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860080678018_390uF
*******
.subckt 860080678019_470uF 1 2
Rser 1 3 0.0232717629338
Lser 2 4 7.313361584E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446809
.ends 860080678019_470uF
*******
.subckt 860080678020_560uF 1 2
Rser 1 3 0.041
Lser 2 4 1.3609256919E-08
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860080678020_560uF
*******
.subckt 860080678021_680uF 1 2
Rser 1 3 0.0199418978859
Lser 2 4 9.773831723E-09
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860080678021_680uF
*******
.subckt 860080678022_820uF 1 2
Rser 1 3 0.0194737704962
Lser 2 4 8.841936425E-09
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860080678022_820uF
*******
.subckt 860080680023_820uF 1 2
Rser 1 3 0.06305
Lser 2 4 1.7911395035E-08
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860080680023_820uF
*******
.subckt 860080680024_1mF 1 2
Rser 1 3 0.0179196008479
Lser 2 4 1.483227424E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 860080680024_1mF
*******
.subckt 860080772001_10uF 1 2
Rser 1 3 0.59
Lser 2 4 0.0000000015
C1 3 4 0.00001
Rpar 3 4 10000000
.ends 860080772001_10uF
*******
.subckt 860080773002_15uF 1 2
Rser 1 3 0.460474259707
Lser 2 4 4.232300922E-09
C1 3 4 0.000015
Rpar 3 4 6666666.66666667
.ends 860080773002_15uF
*******
.subckt 860080773003_18uF 1 2
Rser 1 3 0.32
Lser 2 4 0.0000000028
C1 3 4 0.000018
Rpar 3 4 5555555.55555556
.ends 860080773003_18uF
*******
.subckt 860080773004_22uF 1 2
Rser 1 3 0.339650695071
Lser 2 4 5.189611943E-09
C1 3 4 0.000022
Rpar 3 4 4545454.54545455
.ends 860080773004_22uF
*******
.subckt 860080773005_27uF 1 2
Rser 1 3 0.275709639438
Lser 2 4 3.041167971E-09
C1 3 4 0.000027
Rpar 3 4 3703703.7037037
.ends 860080773005_27uF
*******
.subckt 860080773006_33uF 1 2
Rser 1 3 0.255
Lser 2 4 0.0000000022
C1 3 4 0.000033
Rpar 3 4 3030303.03030303
.ends 860080773006_33uF
*******
.subckt 860080774007_39uF 1 2
Rser 1 3 0.178024439466
Lser 2 4 3.606297262E-09
C1 3 4 0.000039
Rpar 3 4 2564102.56410256
.ends 860080774007_39uF
*******
.subckt 860080774008_47uF 1 2
Rser 1 3 0.147513450046
Lser 2 4 3.965630262E-09
C1 3 4 0.000047
Rpar 3 4 2127659.57446809
.ends 860080774008_47uF
*******
.subckt 860080774009_56uF 1 2
Rser 1 3 0.145
Lser 2 4 0.000000006
C1 3 4 0.000056
Rpar 3 4 1785714.28571429
.ends 860080774009_56uF
*******
.subckt 860080774011_82uF 1 2
Rser 1 3 0.108954873844
Lser 2 4 4.837072923E-09
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860080774011_82uF
*******
.subckt 860080774014_120uF 1 2
Rser 1 3 0.067
Lser 2 4 0.000000007
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860080774014_120uF
*******
.subckt 860080775010_68uF 1 2
Rser 1 3 0.104
Lser 2 4 0.0000000105
C1 3 4 0.000068
Rpar 3 4 1470588.23529412
.ends 860080775010_68uF
*******
.subckt 860080775012_82uF 1 2
Rser 1 3 0.102
Lser 2 4 0.000000009
C1 3 4 0.000082
Rpar 3 4 1219512.19512195
.ends 860080775012_82uF
*******
.subckt 860080775013_100uF 1 2
Rser 1 3 0.100694636813
Lser 2 4 6.447602557E-09
C1 3 4 0.0001
Rpar 3 4 1000000
.ends 860080775013_100uF
*******
.subckt 860080775015_120uF 1 2
Rser 1 3 0.063
Lser 2 4 0.000000007
C1 3 4 0.00012
Rpar 3 4 833333.333333333
.ends 860080775015_120uF
*******
.subckt 860080775016_150uF 1 2
Rser 1 3 0.0791127723048
Lser 2 4 5.611515385E-09
C1 3 4 0.00015
Rpar 3 4 666666.666666667
.ends 860080775016_150uF
*******
.subckt 860080775017_180uF 1 2
Rser 1 3 0.052
Lser 2 4 0.00000001
C1 3 4 0.00018
Rpar 3 4 555555.555555556
.ends 860080775017_180uF
*******
.subckt 860080775018_220uF 1 2
Rser 1 3 0.046
Lser 2 4 0.000000009
C1 3 4 0.00022
Rpar 3 4 454545.454545455
.ends 860080775018_220uF
*******
.subckt 860080775020_330uF 1 2
Rser 1 3 0.0349674626353
Lser 2 4 6.697038625E-09
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080775020_330uF
*******
.subckt 860080778019_270uF 1 2
Rser 1 3 0.0445840995239
Lser 2 4 7.065981861E-09
C1 3 4 0.00027
Rpar 3 4 370370.37037037
.ends 860080778019_270uF
*******
.subckt 860080778021_330uF 1 2
Rser 1 3 0.0340579786939
Lser 2 4 0.000000009400476
C1 3 4 0.00033
Rpar 3 4 303030.303030303
.ends 860080778021_330uF
*******
.subckt 860080778022_390uF 1 2
Rser 1 3 0.0344308769361
Lser 2 4 8.956678893E-09
C1 3 4 0.00039
Rpar 3 4 256410.256410256
.ends 860080778022_390uF
*******
.subckt 860080778023_470uF 1 2
Rser 1 3 0.027156947761
Lser 2 4 8.841934971E-09
C1 3 4 0.00047
Rpar 3 4 212765.957446808
.ends 860080778023_470uF
*******
.subckt 860080780024_470uF 1 2
Rser 1 3 0.0292280789895
Lser 2 4 1.2533114458E-08
C1 3 4 0.00047
Rpar 3 4 212765.957446808
.ends 860080780024_470uF
*******
.subckt 860080780025_560uF 1 2
Rser 1 3 0.0286670439432
Lser 2 4 1.5054867145E-08
C1 3 4 0.00056
Rpar 3 4 178571.428571429
.ends 860080780025_560uF
*******
.subckt 860080780026_680uF 1 2
Rser 1 3 0.0253058048495
Lser 2 4 1.5835711914E-08
C1 3 4 0.00068
Rpar 3 4 147058.823529412
.ends 860080780026_680uF
*******
.subckt 860080780027_820uF 1 2
Rser 1 3 0.0207393465694
Lser 2 4 1.4067758329E-08
C1 3 4 0.00082
Rpar 3 4 121951.219512195
.ends 860080780027_820uF
*******
.subckt 860080780028_1mF 1 2
Rser 1 3 0.0176858108825
Lser 2 4 1.4648292467E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 860080780028_1mF
*******
.subckt 860080781029_1mF 1 2
Rser 1 3 0.0226010170198
Lser 2 4 1.6086029888E-08
C1 3 4 0.001
Rpar 3 4 100000
.ends 860080781029_1mF
*******
.subckt 860080872002_4.7uF 1 2
Rser 1 3 1.3
Lser 2 4 0.000000006
C1 3 4 0.0000047
Rpar 3 4 21276595.7446809
.ends 860080872002_4.7uF
*******
