**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Polymer Capacitors
* Matchcode:             WCAP-PSHP
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 875115150001_220uF 1 2
Rser 1 3 0.00748702469723
Lser 2 4 3.906670607E-09
C1 3 4 0.00022
Rpar 3 4 22727.2727272727
.ends 875115150001_220uF
*******
.subckt 875115150002_270uF 1 2
Rser 1 3 0.010427389814
Lser 2 4 3.929379133E-09
C1 3 4 0.00027
Rpar 3 4 18518.5185185185
.ends 875115150002_270uF
*******
.subckt 875115150003_330uF 1 2
Rser 1 3 0.00915150332731
Lser 2 4 3.726186498E-09
C1 3 4 0.00033
Rpar 3 4 15151.5151515152
.ends 875115150003_330uF
*******
.subckt 875115150004_390uF 1 2
Rser 1 3 0.00714462560492
Lser 2 4 3.842252528E-09
C1 3 4 0.00039
Rpar 3 4 12830.9572301426
.ends 875115150004_390uF
*******
.subckt 875115150005_470uF 1 2
Rser 1 3 0.0131145935317
Lser 2 4 3.844650174E-09
C1 3 4 0.00047
Rpar 3 4 10641.8918918919
.ends 875115150005_470uF
*******
.subckt 875115152006_560uF 1 2
Rser 1 3 0.00881640495169
Lser 2 4 3.812106265E-09
C1 3 4 0.00056
Rpar 3 4 8928.57142857143
.ends 875115152006_560uF
*******
.subckt 875115152007_680uF 1 2
Rser 1 3 0.0133606218464
Lser 2 4 3.827684689E-09
C1 3 4 0.00068
Rpar 3 4 7359.81308411215
.ends 875115152007_680uF
*******
.subckt 875115157010_1.2mF 1 2
Rser 1 3 0.00836577774158
Lser 2 4 5.558365899E-09
C1 3 4 0.0012
Rpar 3 4 5000
.ends 875115157010_1.2mF
*******
.subckt 875115160008_820uF 1 2
Rser 1 3 0.00885045996792
Lser 2 4 4.970322309E-09
C1 3 4 0.00082
Rpar 3 4 6097.56097560976
.ends 875115160008_820uF
*******
.subckt 875115160009_1mF 1 2
Rser 1 3 0.0100331378224
Lser 2 4 5.128608297E-09
C1 3 4 0.001
Rpar 3 4 5000
.ends 875115160009_1mF
*******
.subckt 875115250001_330uF 1 2
Rser 1 3 0.00980553592468
Lser 2 4 3.985487129E-09
C1 3 4 0.00033
Rpar 3 4 15151.5151515152
.ends 875115250001_330uF
*******
.subckt 875115250002_390uF 1 2
Rser 1 3 0.0104900777348
Lser 2 4 3.79968096E-09
C1 3 4 0.00039
Rpar 3 4 12820.5128205128
.ends 875115250002_390uF
*******
.subckt 875115252003_470uF 1 2
Rser 1 3 0.00812051581614
Lser 2 4 3.749982812E-09
C1 3 4 0.00047
Rpar 3 4 10638.2978723404
.ends 875115252003_470uF
*******
.subckt 875115257007_820uF 1 2
Rser 1 3 0.0099813117349
Lser 2 4 5.806855938E-09
C1 3 4 0.00082
Rpar 3 4 6097.56097560976
.ends 875115257007_820uF
*******
.subckt 875115260004_470uF 1 2
Rser 1 3 0.00748648859706
Lser 2 4 5.271611063E-09
C1 3 4 0.00047
Rpar 3 4 10638.2978723404
.ends 875115260004_470uF
*******
.subckt 875115260005_560uF 1 2
Rser 1 3 0.00849483230741
Lser 2 4 5.001273828E-09
C1 3 4 0.00056
Rpar 3 4 8928.57142857143
.ends 875115260005_560uF
*******
.subckt 875115260006_680uF 1 2
Rser 1 3 0.0157281949004
Lser 2 4 4.951514156E-09
C1 3 4 0.00068
Rpar 3 4 7352.94117647059
.ends 875115260006_680uF
*******
.subckt 875115350001_180uF 1 2
Rser 1 3 0.00965391601219
Lser 2 4 3.631797847E-09
C1 3 4 0.00018
Rpar 3 4 55555.5555555556
.ends 875115350001_180uF
*******
.subckt 875115350002_220uF 1 2
Rser 1 3 0.012373298103
Lser 2 4 3.41950618E-09
C1 3 4 0.00022
Rpar 3 4 45454.5454545455
.ends 875115350002_220uF
*******
.subckt 875115352003_270uF 1 2
Rser 1 3 0.01
Lser 2 4 0.0000000025
C1 3 4 0.00027
Rpar 3 4 37037.037037037
.ends 875115352003_270uF
*******
.subckt 875115357006_470uF 1 2
Rser 1 3 0.009
Lser 2 4 0.000000003
C1 3 4 0.00047
Rpar 3 4 21276.5957446809
.ends 875115357006_470uF
*******
.subckt 875115360004_330uF 1 2
Rser 1 3 0.0095
Lser 2 4 0.000000003
C1 3 4 0.00033
Rpar 3 4 30303.0303030303
.ends 875115360004_330uF
*******
.subckt 875115360005_390uF 1 2
Rser 1 3 0.0121300223251
Lser 2 4 4.898103243E-09
C1 3 4 0.00039
Rpar 3 4 25641.0256410256
.ends 875115360005_390uF
*******
.subckt 875115452001_68uF 1 2
Rser 1 3 0.0096888937805
Lser 2 4 3.949628669E-09
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 875115452001_68uF
*******
.subckt 875115452002_82uF 1 2
Rser 1 3 0.00948079243643
Lser 2 4 3.760824407E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 875115452002_82uF
*******
.subckt 875115452003_100uF 1 2
Rser 1 3 0.0106773254387
Lser 2 4 3.606655524E-09
C1 3 4 0.0001
Rpar 3 4 50000
.ends 875115452003_100uF
*******
.subckt 875115452004_150uF 1 2
Rser 1 3 0.0101700335594
Lser 2 4 3.731093687E-09
C1 3 4 0.00015
Rpar 3 4 33333.3333333333
.ends 875115452004_150uF
*******
.subckt 875115457008_270uF 1 2
Rser 1 3 0.0134808650561
Lser 2 4 5.395335774E-09
C1 3 4 0.00027
Rpar 3 4 18518.5185185185
.ends 875115457008_270uF
*******
.subckt 875115460005_150uF 1 2
Rser 1 3 0.0105935646438
Lser 2 4 4.911148019E-09
C1 3 4 0.00015
Rpar 3 4 33333.3333333333
.ends 875115460005_150uF
*******
.subckt 875115460006_180uF 1 2
Rser 1 3 0.0104518653571
Lser 2 4 5.086484187E-09
C1 3 4 0.00018
Rpar 3 4 27777.7777777778
.ends 875115460006_180uF
*******
.subckt 875115460007_220uF 1 2
Rser 1 3 0.0123447747108
Lser 2 4 4.927962554E-09
C1 3 4 0.00022
Rpar 3 4 22727.2727272727
.ends 875115460007_220uF
*******
.subckt 875115552001_68uF 1 2
Rser 1 3 0.0109015046691
Lser 2 4 4.507783507E-09
C1 3 4 0.000068
Rpar 3 4 73529.4117647059
.ends 875115552001_68uF
*******
.subckt 875115552002_82uF 1 2
Rser 1 3 0.0121681202533
Lser 2 4 5.044201258E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 875115552002_82uF
*******
.subckt 875115557005_150uF 1 2
Rser 1 3 0.01
Lser 2 4 5.183210676E-09
C1 3 4 0.00015
Rpar 3 4 33333.3333333333
.ends 875115557005_150uF
*******
.subckt 875115560003_82uF 1 2
Rser 1 3 0.0104243659514
Lser 2 4 5.075291278E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 875115560003_82uF
*******
.subckt 875115560004_100uF 1 2
Rser 1 3 0.0152404870351
Lser 2 4 6.917826409E-09
C1 3 4 0.0001
Rpar 3 4 50000
.ends 875115560004_100uF
*******
.subckt 875115644009_10uF 1 2
Rser 1 3 0.0277297144424
Lser 2 4 2.925731677E-09
C1 3 4 0.00001
Rpar 3 4 58333.3333333333
.ends 875115644009_10uF
*******
.subckt 875115645010_18uF 1 2
Rser 1 3 0.0226811776198
Lser 2 4 3.213299001E-09
C1 3 4 0.000018
Rpar 3 4 58333.3333333333
.ends 875115645010_18uF
*******
.subckt 875115645012_27uF 1 2
Rser 1 3 0.0128005348336
Lser 2 4 2.99640433E-09
C1 3 4 0.000027
Rpar 3 4 58333.3333333333
.ends 875115645012_27uF
*******
.subckt 875115650005_56uF 1 2
Rser 1 3 0.015692292502
Lser 2 4 3.612146676E-09
C1 3 4 0.000056
Rpar 3 4 89285.7142857143
.ends 875115650005_56uF
*******
.subckt 875115652006_82uF 1 2
Rser 1 3 0.0100333339049
Lser 2 4 3.590620949E-09
C1 3 4 0.000082
Rpar 3 4 60975.6097560976
.ends 875115652006_82uF
*******
.subckt 875115652007_100uF 1 2
Rser 1 3 0.0123868521922
Lser 2 4 5.290895138E-09
C1 3 4 0.0001
Rpar 3 4 50000
.ends 875115652007_100uF
*******
.subckt 875115652014_39uF 1 2
Rser 1 3 0.00951131779855
Lser 2 4 3.6772035E-09
C1 3 4 0.000039
Rpar 3 4 58333.3333333333
.ends 875115652014_39uF
*******
.subckt 875115655003_100uF 1 2
Rser 1 3 0.0103
Lser 2 4 0.000000003
C1 3 4 0.0001
Rpar 3 4 869565.217391304
.ends 875115655003_100uF
*******
.subckt 875115655011_22uF 1 2
Rser 1 3 0.0098510988911
Lser 2 4 3.762918893E-09
C1 3 4 0.000022
Rpar 3 4 58333.3333333333
.ends 875115655011_22uF
*******
.subckt 875115655013_33uF 1 2
Rser 1 3 0.00856635233666
Lser 2 4 3.794752483E-09
C1 3 4 0.000033
Rpar 3 4 58333.3333333333
.ends 875115655013_33uF
*******
.subckt 875115655015_56uF 1 2
Rser 1 3 0.0147353075036
Lser 2 4 4.422802993E-09
C1 3 4 0.000056
Rpar 3 4 58333.3333333333
.ends 875115655015_56uF
*******
.subckt 875115657008_120uF 1 2
Rser 1 3 0.0125
Lser 2 4 0.0000000035
C1 3 4 0.00012
Rpar 3 4 41666.6666666667
.ends 875115657008_120uF
*******
.subckt 875115657016_68uF 1 2
Rser 1 3 0.0158804620822
Lser 2 4 5.27053711E-09
C1 3 4 0.000068
Rpar 3 4 58333.3333333333
.ends 875115657016_68uF
*******
.subckt 875115752001_10uF 1 2
Rser 1 3 0.0184012426141
Lser 2 4 5.873354868E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 875115752001_10uF
*******
.subckt 875115852001_10uF 1 2
Rser 1 3 0.0135161211353
Lser 2 4 3.816799008E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 875115852001_10uF
*******
.subckt 875115952001_6.8uF 1 2
Rser 1 3 0.0130576451685
Lser 2 4 3.622186698E-09
C1 3 4 0.0000068
Rpar 3 4 735294.117647059
.ends 875115952001_6.8uF
*******
.subckt 875115957002_12uF 1 2
Rser 1 3 0.0111015775206
Lser 2 4 5.473953262E-09
C1 3 4 0.000012
Rpar 3 4 416666.666666667
.ends 875115957002_12uF
*******
.subckt 875116152001_10uF 1 2
Rser 1 3 0.0149368625192
Lser 2 4 3.730988198E-09
C1 3 4 0.00001
Rpar 3 4 500000
.ends 875116152001_10uF
*******
.subckt 875116157002_15uF 1 2
Rser 1 3 0.0143108149395
Lser 2 4 7.982938621E-09
C1 3 4 0.000015
Rpar 3 4 333333.333333333
.ends 875116157002_15uF
*******
