**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Power Inductor (High Voltage)
* Matchcode:              WE-PD2 HV
* Library Type:           spice
* Version:                rev
* Created/modified by:    Ella
* Date and Time:          7/12/2024
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
.subckt 7850_768775256_560u 1 2
Rp 1 2 135746.824
Cp 1 2 6.3060499p
Rs 1 N3 1.77
L1 N3 2 560u
.ends 7850_768775256_560u
*******
.subckt 7850_768775268_680u 1 2
Rp 1 2 178434.66
Cp 1 2 4.9616929p
Rs 1 N3 2.04
L1 N3 2 680u
.ends 7850_768775268_680u
*******
.subckt 7850_768775282_820u 1 2
Rp 1 2 150782.94
Cp 1 2 4.8144231p
Rs 1 N3 2.35
L1 N3 2 820u
.ends 7850_768775282_820u
*******
.subckt 7850_76877530_1000u 1 2
Rp 1 2 169624.66
Cp 1 2 4.74802404p
Rs 1 N3 2.78
L1 N3 2 1000u
.ends 7850_76877530_1000u
*******
.subckt 7850_768775312_1200u 1 2
Rp 1 2 228952.86
Cp 1 2 5.1586188p
Rs 1 N3 3.77
L1 N3 2 1200u
.ends 7850_768775312_1200u
*******
.subckt 7850_768775322_2200u 1 2
Rp 1 2 225324.09
Cp 1 2 5.2462005p
Rs 1 N3 6
L1 N3 2 2200u
.ends 7850_768775322_2200u
*******
.subckt 1054_76877630_1000u 1 2
Rp 1 2 230366
Cp 1 2 4.954p
Rs 1 N3 2.2
L1 N3 2 1000u
.ends 1054_76877630_1000u
*******
.subckt 1054_768776312_1200u 1 2
Rp 1 2 165813.51
Cp 1 2 5.4492682p
Rs 1 N3 2.48
L1 N3 2 1200u
.ends 1054_768776312_1200u
*******
.subckt 1054_768776322_2200u 1 2
Rp 1 2 275669.169519
Cp 1 2 5.33990012326p
Rs 1 N3 4.4
L1 N3 2 2200u
.ends 1054_768776322_2200u
*******
