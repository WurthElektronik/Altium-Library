**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 Aluminum Polymer Capacitors
* Matchcode:             WCAP-PSLP
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         6/1/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 875105142001_47uF 1 2
Rser 1 3 0.0146178023095
Lser 2 4 3.503849781E-09
C1 3 4 0.000047
Rpar 3 4 21000
.ends 875105142001_47uF
*******
.subckt 875105142002_56uF 1 2
Rser 1 3 0.0159256096044
Lser 2 4 2.761083171E-09
C1 3 4 0.000056
Rpar 3 4 21000
.ends 875105142002_56uF
*******
.subckt 875105142003_68uF 1 2
Rser 1 3 0.0125948257859
Lser 2 4 2.79992293E-09
C1 3 4 0.000068
Rpar 3 4 21000
.ends 875105142003_68uF
*******
.subckt 875105142004_82uF 1 2
Rser 1 3 0.0142038332755
Lser 2 4 2.832972153E-09
C1 3 4 0.000082
Rpar 3 4 21000
.ends 875105142004_82uF
*******
.subckt 875105142005_100uF 1 2
Rser 1 3 0.0101849521435
Lser 2 4 2.730940001E-09
C1 3 4 0.0001
Rpar 3 4 21000
.ends 875105142005_100uF
*******
.subckt 875105142006_150uF 1 2
Rser 1 3 0.0112204509376
Lser 2 4 2.612408389E-09
C1 3 4 0.00015
Rpar 3 4 21000
.ends 875105142006_150uF
*******
.subckt 875105144007_180uF 1 2
Rser 1 3 0.00918784444536
Lser 2 4 2.991114514E-09
C1 3 4 0.00018
Rpar 3 4 21000
.ends 875105144007_180uF
*******
.subckt 875105144008_220uF 1 2
Rser 1 3 0.0119373056532
Lser 2 4 3.001034672E-09
C1 3 4 0.00022
Rpar 3 4 21000
.ends 875105144008_220uF
*******
.subckt 875105144009_270uF 1 2
Rser 1 3 0.0126993981475
Lser 2 4 3.470113431E-09
C1 3 4 0.00027
Rpar 3 4 21000
.ends 875105144009_270uF
*******
.subckt 875105144010_330uF 1 2
Rser 1 3 0.0165611581005
Lser 2 4 3.005418053E-09
C1 3 4 0.00033
Rpar 3 4 21000
.ends 875105144010_330uF
*******
.subckt 875105145011_390uF 1 2
Rser 1 3 0.00950335433369
Lser 2 4 3.23809525E-09
C1 3 4 0.00039
Rpar 3 4 21000
.ends 875105145011_390uF
*******
.subckt 875105240001_10uF 1 2
Rser 1 3 0.018084356216
Lser 2 4 2.335490858E-09
C1 3 4 0.00001
Rpar 3 4 33333.3333333333
.ends 875105240001_10uF
*******
.subckt 875105240002_15uF 1 2
Rser 1 3 0.0159479420491
Lser 2 4 2.361682514E-09
C1 3 4 0.000015
Rpar 3 4 33333.3333333333
.ends 875105240002_15uF
*******
.subckt 875105240003_22uF 1 2
Rser 1 3 0.0186709974457
Lser 2 4 2.448962924E-09
C1 3 4 0.000022
Rpar 3 4 33333.3333333333
.ends 875105240003_22uF
*******
.subckt 875105242004_33uF 1 2
Rser 1 3 0.0219163226283
Lser 2 4 2.859600019E-09
C1 3 4 0.000033
Rpar 3 4 33333.3333333333
.ends 875105242004_33uF
*******
.subckt 875105242005_39uF 1 2
Rser 1 3 0.0146268318602
Lser 2 4 2.546390513E-09
C1 3 4 0.000039
Rpar 3 4 33333.3333333333
.ends 875105242005_39uF
*******
.subckt 875105242006_47uF 1 2
Rser 1 3 0.023226581579
Lser 2 4 3.137650187E-09
C1 3 4 0.000047
Rpar 3 4 33333.3333333333
.ends 875105242006_47uF
*******
.subckt 875105242007_56uF 1 2
Rser 1 3 0.012296122735
Lser 2 4 2.638679056E-09
C1 3 4 0.000056
Rpar 3 4 33333.3333333333
.ends 875105242007_56uF
*******
.subckt 875105242008_68uF 1 2
Rser 1 3 0.0115729421122
Lser 2 4 2.678751815E-09
C1 3 4 0.000068
Rpar 3 4 33333.3333333333
.ends 875105242008_68uF
*******
.subckt 875105242009_82uF 1 2
Rser 1 3 0.01766
Lser 2 4 2.44417180868638E-09
C1 3 4 0.000082
Rpar 3 4 33333.3333333333
.ends 875105242009_82uF
*******
.subckt 875105242010_100uF 1 2
Rser 1 3 0.0124059822172
Lser 2 4 2.715206427E-09
C1 3 4 0.0001
Rpar 3 4 33333.3333333333
.ends 875105242010_100uF
*******
.subckt 875105244011_150uF 1 2
Rser 1 3 0.0106479827332
Lser 2 4 2.86665223E-09
C1 3 4 0.00015
Rpar 3 4 33333.3333333333
.ends 875105244011_150uF
*******
.subckt 875105244012_180uF 1 2
Rser 1 3 0.0242796156982
Lser 2 4 3.298908307E-09
C1 3 4 0.00018
Rpar 3 4 33333.3333333333
.ends 875105244012_180uF
*******
.subckt 875105244013_220uF 1 2
Rser 1 3 0.0114523311763
Lser 2 4 2.845376354E-09
C1 3 4 0.00022
Rpar 3 4 33333.3333333333
.ends 875105244013_220uF
*******
.subckt 875105245014_270uF 1 2
Rser 1 3 0.0108531159206
Lser 2 4 3.321753848E-09
C1 3 4 0.00027
Rpar 3 4 33333.3333333333
.ends 875105245014_270uF
*******
.subckt 875105245015_330uF 1 2
Rser 1 3 0.0113192832289
Lser 2 4 3.374454181E-09
C1 3 4 0.00033
Rpar 3 4 33333.3333333333
.ends 875105245015_330uF
*******
.subckt 875105344006_47uF 1 2
Rser 1 3 0.0211025530363
Lser 2 4 3.090667045E-09
C1 3 4 0.000047
Rpar 3 4 40000
.ends 875105344006_47uF
*******
.subckt 875105344007_56uF 1 2
Rser 1 3 0.0113095080484
Lser 2 4 3.032659201E-09
C1 3 4 0.000056
Rpar 3 4 40000
.ends 875105344007_56uF
*******
.subckt 875105344008_68uF 1 2
Rser 1 3 0.0237335503052
Lser 2 4 3.297798943E-09
C1 3 4 0.000068
Rpar 3 4 40000
.ends 875105344008_68uF
*******
.subckt 875105344009_82uF 1 2
Rser 1 3 0.0158485046548
Lser 2 4 2.897198281E-09
C1 3 4 0.000082
Rpar 3 4 40000
.ends 875105344009_82uF
*******
.subckt 875105344010_100uF 1 2
Rser 1 3 0.0163097755095
Lser 2 4 3.124563497E-09
C1 3 4 0.0001
Rpar 3 4 40000
.ends 875105344010_100uF
*******
.subckt 875105345011_150uF 1 2
Rser 1 3 0.0119350945534
Lser 2 4 3.098422093E-09
C1 3 4 0.00015
Rpar 3 4 40000
.ends 875105345011_150uF
*******
.subckt 875105359001_10uF 1 2
Rser 1 3 0.0191074985904
Lser 2 4 2.619590372E-09
C1 3 4 0.00001
Rpar 3 4 40000
.ends 875105359001_10uF
*******
.subckt 875105359002_15uF 1 2
Rser 1 3 0.0165014517982
Lser 2 4 2.538922307E-09
C1 3 4 0.000015
Rpar 3 4 40000
.ends 875105359002_15uF
*******
.subckt 875105359003_22uF 1 2
Rser 1 3 0.0169707022759
Lser 2 4 2.466059541E-09
C1 3 4 0.000022
Rpar 3 4 40000
.ends 875105359003_22uF
*******
.subckt 875105359004_33uF 1 2
Rser 1 3 0.0165101149951
Lser 2 4 2.54913326E-09
C1 3 4 0.000033
Rpar 3 4 40000
.ends 875105359004_33uF
*******
.subckt 875105359005_39uF 1 2
Rser 1 3 0.0191964937563
Lser 2 4 2.639803204E-09
C1 3 4 0.000039
Rpar 3 4 40000
.ends 875105359005_39uF
*******
.subckt 875105444001_10uF 1 2
Rser 1 3 0.0276978442436
Lser 2 4 3.245492716E-09
C1 3 4 0.00001
Rpar 3 4 33333.3333333333
.ends 875105444001_10uF
*******
.subckt 875105444002_15uF 1 2
Rser 1 3 0.0146050544329
Lser 2 4 3.22977463E-09
C1 3 4 0.000015
Rpar 3 4 33333.3333333333
.ends 875105444002_15uF
*******
.subckt 875105444003_22uF 1 2
Rser 1 3 0.0191932128155
Lser 2 4 2.995436701E-09
C1 3 4 0.000022
Rpar 3 4 33333.3333333333
.ends 875105444003_22uF
*******
.subckt 875105444004_33uF 1 2
Rser 1 3 0.0167661846845
Lser 2 4 3.015220567E-09
C1 3 4 0.000033
Rpar 3 4 33333.3333333333
.ends 875105444004_33uF
*******
.subckt 875105445005_39uF 1 2
Rser 1 3 0.0107445722067
Lser 2 4 3.258401177E-09
C1 3 4 0.000039
Rpar 3 4 33333.3333333333
.ends 875105445005_39uF
*******
.subckt 875105445006_47uF 1 2
Rser 1 3 0.0115087958692
Lser 2 4 3.235775785E-09
C1 3 4 0.000047
Rpar 3 4 33333.3333333333
.ends 875105445006_47uF
*******
.subckt 875105445007_56uF 1 2
Rser 1 3 0.0187928809704
Lser 2 4 3.508500669E-09
C1 3 4 0.000056
Rpar 3 4 33333.3333333333
.ends 875105445007_56uF
*******
.subckt 875105544001_10uF 1 2
Rser 1 3 0.0204482140593
Lser 2 4 3.010157832E-09
C1 3 4 0.00001
Rpar 3 4 41666.6666666667
.ends 875105544001_10uF
*******
.subckt 875105544002_15uF 1 2
Rser 1 3 0.0184587224254
Lser 2 4 2.834629347E-09
C1 3 4 0.000015
Rpar 3 4 41666.6666666667
.ends 875105544002_15uF
*******
.subckt 875105544003_22uF 1 2
Rser 1 3 0.0196880023174
Lser 2 4 2.964470061E-09
C1 3 4 0.000022
Rpar 3 4 41666.6666666667
.ends 875105544003_22uF
*******
.subckt 875105545004_33uF 1 2
Rser 1 3 0.0182318807924
Lser 2 4 4.406523353E-09
C1 3 4 0.000033
Rpar 3 4 41666.6666666667
.ends 875105545004_33uF
*******
.subckt 875105545005_39uF 1 2
Rser 1 3 0.0149915964408
Lser 2 4 3.50316725E-09
C1 3 4 0.000039
Rpar 3 4 41666.6666666667
.ends 875105545005_39uF
*******
.subckt 875105644004_18uF 1 2
Rser 1 3 0.0296469307671
Lser 2 4 3.763764556E-09
C1 3 4 0.000018
Rpar 3 4 58333.3333333333
.ends 875105644004_18uF
*******
.subckt 875105645005_47uF 1 2
Rser 1 3 0.0139460850391
Lser 2 4 3.258713889E-09
C1 3 4 0.000047
Rpar 3 4 58333.3333333333
.ends 875105645005_47uF
*******
.subckt 875105744001_8.2uF 1 2
Rser 1 3 0.0377957322814
Lser 2 4 2.943717326E-09
C1 3 4 0.0000082
Rpar 3 4 83333.3333333333
.ends 875105744001_8.2uF
*******
.subckt 875105744002_12uF 1 2
Rser 1 3 0.0425392751929
Lser 2 4 4.325234269E-09
C1 3 4 0.000012
Rpar 3 4 83333.3333333333
.ends 875105744002_12uF
*******
.subckt 875105744003_15uF 1 2
Rser 1 3 0.0290464276906
Lser 2 4 4.622002884E-09
C1 3 4 0.000015
Rpar 3 4 83333.3333333333
.ends 875105744003_15uF
*******
.subckt 875105844001_5.6uF 1 2
Rser 1 3 0.0325200282212
Lser 2 4 3.177951647E-09
C1 3 4 0.0000056
Rpar 3 4 105000
.ends 875105844001_5.6uF
*******
.subckt 875105844002_8.2uF 1 2
Rser 1 3 0.0363051600961
Lser 2 4 2.812410146E-09
C1 3 4 0.0000082
Rpar 3 4 105000
.ends 875105844002_8.2uF
*******
.subckt 875105945001_4.7uF 1 2
Rser 1 3 0.0100333339049
Lser 2 4 3.590620949E-09
C1 3 4 0.0000047
Rpar 3 4 166666.666666667
.ends 875105945001_4.7uF
*******
