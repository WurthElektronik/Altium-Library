**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Infrared Ceramic Waterclear
* Matchcode:              WL-SIMW
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-03-01
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 3535_15435385A9050  1  2
D1 1 2 SIMW
.MODEL SIMW D
+ IS=10.000E-21
+ N=1.2042
+ RS=.62459
+ IKF=.16435
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt 3535_15435385AA350  1  2
D1 1 2 SIMW
.MODEL SIMW D
+ IS=44.425E-21
+ N=1.2686
+ RS=.84728
+ IKF=249.76
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt  3535_15435394A9050  1  2
D1 1 2 SIMW
.MODEL SIMW D
+ IS=10.000E-21
+ N=1.0843
+ RS=.51194
+ IKF=.27452
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******
.subckt  3535_15435394AA350  1  2
D1 1 2 SIMW
.MODEL SIMW D
+ IS=10.000E-21
+ N=1.0916
+ RS=.54324
+ IKF=.20186
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=5
+ IBV=10.00E-6
+ TT=5.0000E-9
.ends
******