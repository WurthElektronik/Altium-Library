**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  SMT Power Inductor
* Matchcode:              WE-PD3
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-06-10
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt TypeL_74454010_10u 1 2
Rp 1 2 14450
Cp 1 2 4.55p
Rs 1 N3 0.048
L1 N3 2 10u
.ends TypeL_74454010_10u
*******
.subckt TypeL_7445402_2.2u 1 2
Rp 1 2 3900
Cp 1 2 1.7p
Rs 1 N3 0.023
L1 N3 2 2.2u
.ends TypeL_7445402_2.2u
*******
.subckt TypeL_7445403_3u 1 2
Rp 1 2 5250
Cp 1 2 1.85p
Rs 1 N3 0.026
L1 N3 2 3u
.ends TypeL_7445403_3u
*******
.subckt TypeL_7445404_4.7u 1 2
Rp 1 2 8650
Cp 1 2 2.1p
Rs 1 N3 0.034
L1 N3 2 4.7u
.ends TypeL_7445404_4.7u
*******
.subckt TypeL_74454068_7u 1 2
Rp 1 2 11100
Cp 1 2 3.7p
Rs 1 N3 0.041
L1 N3 2 7u
.ends TypeL_74454068_7u
*******
.subckt TypeL_74454115_15u 1 2
Rp 1 2 19400
Cp 1 2 4.3p
Rs 1 N3 0.064
L1 N3 2 15u
.ends TypeL_74454115_15u
*******
.subckt TypeL_74454122_22u 1 2
Rp 1 2 23300
Cp 1 2 4.5p
Rs 1 N3 0.076
L1 N3 2 22u
.ends TypeL_74454122_22u
*******
.subckt TypeL_74454133_33u 1 2
Rp 1 2 36000
Cp 1 2 6.4p
Rs 1 N3 0.127
L1 N3 2 33u
.ends TypeL_74454133_33u
*******
.subckt TypeL_74454147_47u 1 2
Rp 1 2 51150
Cp 1 2 5.4p
Rs 1 N3 0.158
L1 N3 2 47u
.ends TypeL_74454147_47u
*******
.subckt TypeL_74454168_68u 1 2
Rp 1 2 64300
Cp 1 2 6p
Rs 1 N3 0.285
L1 N3 2 68u
.ends TypeL_74454168_68u
*******
.subckt TypeL_7445420_100u 1 2
Rp 1 2 108850
Cp 1 2 4.7p
Rs 1 N3 0.373
L1 N3 2 100u
.ends TypeL_7445420_100u
*******
.subckt TypeL_74454215_150u 1 2
Rp 1 2 115150
Cp 1 2 5p
Rs 1 N3 0.456
L1 N3 2 150u
.ends TypeL_74454215_150u
*******
.subckt TypeL_74454220_220u 1 2
Rp 1 2 145900
Cp 1 2 5.65p
Rs 1 N3 0.683
L1 N3 2 220u
.ends TypeL_74454220_220u
*******
.subckt TypeL_74454233_330u 1 2
Rp 1 2 160950
Cp 1 2 7.4p
Rs 1 N3 1.044
L1 N3 2 330u
.ends TypeL_74454233_330u
*******
.subckt TypeL_74454239_390u 1 2
Rp 1 2 168150
Cp 1 2 5.7p
Rs 1 N3 1.175
L1 N3 2 390u
.ends TypeL_74454239_390u
*******
.subckt TypeL_74454247_470u 1 2
Rp 1 2 204750
Cp 1 2 5.4p
Rs 1 N3 1.35
L1 N3 2 470u
.ends TypeL_74454247_470u
*******
.subckt TypeL_74454268_680u 1 2
Rp 1 2 220700
Cp 1 2 6.4p
Rs 1 N3 1.94
L1 N3 2 680u
.ends TypeL_74454268_680u
*******
.subckt TypeL_7445430_1m 1 2
Rp 1 2 282800
Cp 1 2 5.3p
Rs 1 N3 2.75
L1 N3 2 1000u
.ends TypeL_7445430_1m
*******
.subckt TypeM_7445301_1.5u 1 2
Rp 1 2 3125
Cp 1 2 1.95p
Rs 1 N3 0.029
L1 N3 2 1.5u
.ends TypeM_7445301_1.5u
*******
.subckt TypeM_74453010_10u 1 2
Rp 1 2 10150
Cp 1 2 3.6p
Rs 1 N3 0.117
L1 N3 2 10u
.ends TypeM_74453010_10u
*******
.subckt TypeM_7445302_2.2u 1 2
Rp 1 2 4950
Cp 1 2 2.2p
Rs 1 N3 0.037
L1 N3 2 2.2u
.ends TypeM_7445302_2.2u
*******
.subckt TypeM_7445303_3.9u 1 2
Rp 1 2 8500
Cp 1 2 2.8p
Rs 1 N3 0.058
L1 N3 2 3.9u
.ends TypeM_7445303_3.9u
*******
.subckt TypeM_74453031_3.3u 1 2
Rp 1 2 8195
Cp 1 2 2.6p
Rs 1 N3 0.052
L1 N3 2 3.3u
.ends TypeM_74453031_3.3u
*******
.subckt TypeM_7445304_4.7u 1 2
Rp 1 2 8800
Cp 1 2 2.9p
Rs 1 N3 0.065
L1 N3 2 4.7u
.ends TypeM_7445304_4.7u
*******
.subckt TypeM_7445306_6.8u 1 2
Rp 1 2 8550
Cp 1 2 3.1p
Rs 1 N3 0.064
L1 N3 2 6.8u
.ends TypeM_7445306_6.8u
*******
.subckt TypeM_74453112_12u 1 2
Rp 1 2 13350
Cp 1 2 3.3p
Rs 1 N3 0.16
L1 N3 2 12u
.ends TypeM_74453112_12u
*******
.subckt TypeM_74453115_15u 1 2
Rp 1 2 15750
Cp 1 2 3.5p
Rs 1 N3 0.17
L1 N3 2 15u
.ends TypeM_74453115_15u
*******
.subckt TypeM_74453122_22u 1 2
Rp 1 2 17450
Cp 1 2 3.4p
Rs 1 N3 0.248
L1 N3 2 22u
.ends TypeM_74453122_22u
*******
.subckt TypeM_74453133_33u 1 2
Rp 1 2 25840
Cp 1 2 3.3p
Rs 1 N3 0.371
L1 N3 2 33u
.ends TypeM_74453133_33u
*******
.subckt TypeM_74453147_47u 1 2
Rp 1 2 31850
Cp 1 2 3.2p
Rs 1 N3 0.481
L1 N3 2 47u
.ends TypeM_74453147_47u
*******
.subckt TypeM_74453156_56u 1 2
Rp 1 2 36900
Cp 1 2 4p
Rs 1 N3 0.552
L1 N3 2 56u
.ends TypeM_74453156_56u
*******
.subckt TypeM_74453168_68u 1 2
Rp 1 2 38700
Cp 1 2 4p
Rs 1 N3 0.62
L1 N3 2 68u
.ends TypeM_74453168_68u
*******
.subckt TypeM_74453182_82u 1 2
Rp 1 2 46800
Cp 1 2 3.8p
Rs 1 N3 1.03
L1 N3 2 82u
.ends TypeM_74453182_82u
*******
.subckt TypeM_7445320_100u 1 2
Rp 1 2 53650
Cp 1 2 4.3p
Rs 1 N3 1.164
L1 N3 2 100u
.ends TypeM_7445320_100u
*******
.subckt TypeS_7445101_1u 1 2
Rp 1 2 380
Cp 1 2 0.635p
Rs 1 N3 0.014
L1 N3 2 1u
.ends TypeS_7445101_1u
*******
.subckt TypeS_74451015_1.5u 1 2
Rp 1 2 600
Cp 1 2 0.985p
Rs 1 N3 0.018
L1 N3 2 1.5u
.ends TypeS_74451015_1.5u
*******
.subckt TypeS_74451022_2.2u 1 2
Rp 1 2 715
Cp 1 2 1.14p
Rs 1 N3 0.021
L1 N3 2 2.2u
.ends TypeS_74451022_2.2u
*******
.subckt TypeS_74451033_3.3u 1 2
Rp 1 2 1230
Cp 1 2 1.23p
Rs 1 N3 0.025
L1 N3 2 3.3u
.ends TypeS_74451033_3.3u
*******
.subckt TypeS_74451039_4.3u 1 2
Rp 1 2 1570
Cp 1 2 1.53p
Rs 1 N3 0.04
L1 N3 2 4.3u
.ends TypeS_74451039_4.3u
*******
.subckt TypeS_74451047_4.7u 1 2
Rp 1 2 1880
Cp 1 2 2.05p
Rs 1 N3 0.045
L1 N3 2 4.7u
.ends TypeS_74451047_4.7u
*******
.subckt TypeS_74451068_6.8u 1 2
Rp 1 2 2230
Cp 1 2 2.277p
Rs 1 N3 0.055
L1 N3 2 6.8u
.ends TypeS_74451068_6.8u
*******
.subckt TypeS_7445110_10u 1 2
Rp 1 2 2830
Cp 1 2 2.8p
Rs 1 N3 0.056
L1 N3 2 10u
.ends TypeS_7445110_10u
*******
.subckt TypeS_74451115_15u 1 2
Rp 1 2 3200
Cp 1 2 3.13p
Rs 1 N3 0.075
L1 N3 2 15u
.ends TypeS_74451115_15u
*******
.subckt TypeS_74451122_22u 1 2
Rp 1 2 7400
Cp 1 2 3.3p
Rs 1 N3 0.09
L1 N3 2 22u
.ends TypeS_74451122_22u
*******
.subckt TypeS_74451133_33u 1 2
Rp 1 2 7800
Cp 1 2 3.6p
Rs 1 N3 0.114
L1 N3 2 33u
.ends TypeS_74451133_33u
*******
.subckt TypeS_74451147_47u 1 2
Rp 1 2 9000
Cp 1 2 3.9p
Rs 1 N3 0.16
L1 N3 2 47u
.ends TypeS_74451147_47u
*******
.subckt TypeS_74451168_68u 1 2
Rp 1 2 10600
Cp 1 2 4.3p
Rs 1 N3 0.221
L1 N3 2 68u
.ends TypeS_74451168_68u
*******
.subckt TypeS_7445120_100u 1 2
Rp 1 2 15200
Cp 1 2 3.74p
Rs 1 N3 0.393
L1 N3 2 100u
.ends TypeS_7445120_100u
*******
.subckt TypeS_74451215_150u 1 2
Rp 1 2 14000
Cp 1 2 4.7p
Rs 1 N3 0.41
L1 N3 2 150u
.ends TypeS_74451215_150u
*******
.subckt TypeS_74451222_220u 1 2
Rp 1 2 17000
Cp 1 2 5p
Rs 1 N3 0.58
L1 N3 2 220u
.ends TypeS_74451222_220u
*******
.subckt TypeS_74451233_330u 1 2
Rp 1 2 29000
Cp 1 2 5.3p
Rs 1 N3 1
L1 N3 2 330u
.ends TypeS_74451233_330u
*******
.subckt TypeS_74451247_470u 1 2
Rp 1 2 42000
Cp 1 2 6.5p
Rs 1 N3 1.7
L1 N3 2 470u
.ends TypeS_74451247_470u
*******
.subckt TypeX_74459010_10u 1 2
Rp 1 2 12100
Cp 1 2 5.35p
Rs 1 N3 0.023
L1 N3 2 10u
.ends TypeX_74459010_10u
*******
.subckt TypeX_74459115_15u 1 2
Rp 1 2 12740
Cp 1 2 6.15p
Rs 1 N3 0.03
L1 N3 2 15u
.ends TypeX_74459115_15u
*******
.subckt TypeX_74459122_22u 1 2
Rp 1 2 21800
Cp 1 2 6.5p
Rs 1 N3 0.048
L1 N3 2 22u
.ends TypeX_74459122_22u
*******
.subckt TypeX_74459133_33u 1 2
Rp 1 2 27850
Cp 1 2 6.6p
Rs 1 N3 0.071
L1 N3 2 33u
.ends TypeX_74459133_33u
*******
.subckt TypeX_74459147_47u 1 2
Rp 1 2 35350
Cp 1 2 8p
Rs 1 N3 0.085
L1 N3 2 47u
.ends TypeX_74459147_47u
*******
.subckt TypeX_74459168_68u 1 2
Rp 1 2 65200
Cp 1 2 7.1p
Rs 1 N3 0.105
L1 N3 2 68u
.ends TypeX_74459168_68u
*******
.subckt TypeX_7445920_100u 1 2
Rp 1 2 90850
Cp 1 2 8.5p
Rs 1 N3 0.151
L1 N3 2 100u
.ends TypeX_7445920_100u
*******
.subckt TypeX_74459215_150u 1 2
Rp 1 2 94350
Cp 1 2 8.9p
Rs 1 N3 0.209
L1 N3 2 150u
.ends TypeX_74459215_150u
*******
.subckt TypeX_74459222_220u 1 2
Rp 1 2 101350
Cp 1 2 10.15p
Rs 1 N3 0.311
L1 N3 2 220u
.ends TypeX_74459222_220u
*******
.subckt TypeX_74459233_330u 1 2
Rp 1 2 115950
Cp 1 2 9.8p
Rs 1 N3 0.457
L1 N3 2 330u
.ends TypeX_74459233_330u
*******
.subckt TypeX_74459247_470u 1 2
Rp 1 2 129600
Cp 1 2 10p
Rs 1 N3 0.661
L1 N3 2 470u
.ends TypeX_74459247_470u
*******
.subckt TypeX_74459268_680u 1 2
Rp 1 2 183950
Cp 1 2 8.6p
Rs 1 N3 1.059
L1 N3 2 680u
.ends TypeX_74459268_680u
*******
.subckt TypeX_7445930_1m 1 2
Rp 1 2 218500
Cp 1 2 9p
Rs 1 N3 1.427
L1 N3 2 1000u
.ends TypeX_7445930_1m
*******
