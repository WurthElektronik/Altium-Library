**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Energy Harvesting Coupled Inductor
* Matchcode:              WE-EHPI 
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-05-25
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 5838_74488540250_25u  1  2  3  4  PARAMS:
+  Cww=7.92p
+  Rp1=1694
+  Cp1=3.793n
+  Lp1=24.543u
+  Rp2=656715
+  Cp2=11.347p
+  Lp2=10.366m
+  RDC1=0.040
+  RDC2=0.2
+  K=0.97899637
C_C1  1  4    {Cww/2}
C_C2  2  3    {Cww/2}
C_C5  2  1    {Cp1}
R_R1  2  N05454    {RDC1}
R_R2  2  1    {Rp1}
L_L1  N05454  1    {Lp1}
L_L2  N05750  4    {Lp2}
C_C6  3  4    {Cp2}
R_R3  3  4    {Rp2}
R_R4  3  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
**************************************************
.subckt 5838_74488540120_13u  1  2  3  4  PARAMS:
+  Cww=6.28p
+  Rp1=550
+  Cp1=17n
+  Lp1=13.01u
+  Rp2=275585
+  Cp2=8.98p
+  Lp2=33.116m
+  RDC1=0.135
+  RDC2=0.09
+  K=0.975605608
C_C1  1  4    {Cww/2}
C_C2  2  3    {Cww/2}
C_C5  2  1    {Cp1}
R_R1  2  N05454    {RDC1}
R_R2  2  1    {Rp1}
L_L1  N05454  1    {Lp1}
L_L2  N05750  4    {Lp2}
C_C6  3  4    {Cp2}
R_R3  3  4    {Rp2}
R_R4  3  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
**************************************************
.subckt 5838_74488540070_7u  1  2  3  4  PARAMS:
+  Cww=6.91p
+  Rp1=280
+  Cp1=70n
+  Lp1=6.8u
+  Rp2=248260
+  Cp2=8.797p
+  Lp2=69.487m
+  RDC1=0.205
+  RDC2=0.085
+  K=0.969535971
C_C1  1  4    {Cww/2}
C_C2  2  3    {Cww/2}
C_C5  2  1    {Cp1}
R_R1  2  N05454    {RDC1}
R_R2  2  1    {Rp1}
L_L1  N05454  1    {Lp1}
L_L2  N05750  4    {Lp2}
C_C6  3  4    {Cp2}
R_R3  3  4    {Rp2}
R_R4  3  N05750    {RDC2}
Kn_K1  L_L1  L_L2      {K}
.ends
******