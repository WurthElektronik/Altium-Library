**************************************************
* Manufacturer:           Wurth Elektronik 
* Kinds:                  Optocoupler Darlington
* Matchcode:              WL-OCDA
* Library Type:           LTspice
* Version:                rev22a
* Created/modified by:    Ella      
* Date and Time:          2022-02-14
* Team:                   eiSos EDA Service  
* Contact:                libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.SUBCKT Series_352_14135214xxx A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.003,
+ (0.12010E-02*EXP(-0.13696E+02*EXP(-0.43553E+04*V(T)))-0.51169E-05)/100,
+ (-0.693889E-17*V(T)+0.119524E-02)/100)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=121.43E-18
+ N=1.4750
+ RS=1.3001
+ IKF=.22024
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9

.model Detector NPN IS=3.64P BF=8000 NF=2 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=200 IKF=20 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_815_14181514xxx A K C E 
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.003,
+ (0.13594E-02/(1+0.70683E+01*EXP(-0.38001E+04*V(T)))-0.17655E-03)/100,
+ (0.254110E-20/V(T)+0.117988E-02)/100)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=22.505E-18
+ N=1.4098
+ RS=.47806
+ IKF=17.001E-3
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9

.model Detector NPN IS=3.64P BF=3500 NF=1.24 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=100 IKF=10 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************
.SUBCKT Series_355_14135514xxx A K C E
D1 A D LED	
VH D K 0 
Hd R 0 VH 1	
Rd R T 10k
Cd T 0 0.02n
Rg B 0 4G
Q1 C B E Detector

G1 C B TABLE
+ {if(V(T)<0.003,
+ (0.15076E-02/(1+0.10831E+02*EXP(-0.35692E+04*V(T)))-0.15409E-03)/100,
+ (-0.254110E-20/V(T)+0.134724E-02)/100)}
+ (0,0.0000000001) (10,10)

.model LED D
+ IS=566.88E-18
+ N=1.5480
+ RS=1.1990
+ CJO=1.0000E-12
+ M=.3333
+ VJ=.75
+ BV=6
+ IBV=10.00E-6
+ TT=5.0000E-9

.model Detector NPN IS=3.64P BF=3500 NF=1.265 BR=10 TF=20N TR=350n
+ CJE=5.16P VJE=0.99 MJE=0.2411274 CJC=18P VJC=0.597478 MJC=0.431978
+ ISC=0.207N VAF=300 IKF=200 ISS=0 CJS=7.74p VJS=0.61 MJS=0.31
.ends
***********************