**************************************************
* Manufacturer:          Wurth Elektronik 
* Kinds:                 SMT EMI Suppression Power Ferrite
* Matchcode:             WE-PF
* Library Type:          LTspice
* Version:               rev22a
* Created/modified by:   Ella
* Date and Time:         5/30/2022
* Team:                  eiSos EDA Service  
* Contact:               libraries@we-online.com
**************************************************
* Copyright(C) 2022 Würth Elektronik eiSos GmbH & Co. KG
* All Rights Reserved.
**************************************************
* Disclaimer: While Würth Elektronik eiSos has made every reasonable effort to ensure the accuracy
* of the simulation models provided, Würth Elektronik eiSos does not guarantee the exemption of error on
* the simulation models, nor does Würth Elektronik eiSos guarantee that the simulation model is current.
* Würth Elektronik eiSos reserves the right to make any adjustments at any time without notice.
* Würth Elektronik eiSos expressly disclaims all implied warranties regarding this simulation model.
**************************************************
.subckt 1280_742792901_1180ohm 1 2
Rp 1 2 1830
Cp 1 2 4.026p
Rs 1 N3 0.009
L1 N3 2 0.796071u
.ends 1280_742792901_1180ohm
*******
.subckt 1280_742792902_565ohm 1 2
Rp 1 2 3964
Cp 1 2 2.41p
Rs 1 N3 0.012
L1 N3 2 2.187u
.ends 1280_742792902_565ohm
*******
.subckt 1280_742792903_340ohm 1 2
Rp 1 2 4310
Cp 1 2 6.73p
Rs 1 N3 0.009
L1 N3 2 2.801u
.ends 1280_742792903_340ohm
*******
.subckt 1280_742792904_300ohm 1 2
Rp 1 2 4621
Cp 1 2 8.065p
Rs 1 N3 0.015
L1 N3 2 3.414u
.ends 1280_742792904_300ohm
*******
.subckt 1280_742792906_190ohm 1 2
Rp 1 2 5933
Cp 1 2 13.8p
Rs 1 N3 0.02
L1 N3 2 4.574u
.ends 1280_742792906_190ohm
*******
.subckt 1280_742792907_240ohm 1 2
Rp 1 2 6588
Cp 1 2 10.104p
Rs 1 N3 0.02
L1 N3 2 6.222u
.ends 1280_742792907_240ohm
*******
.subckt 1280_742792910_200ohm 1 2
Rp 1 2 6399
Cp 1 2 4.71p
Rs 1 N3 0.025
L1 N3 2 8.662u
.ends 1280_742792910_200ohm
*******
.subckt 1280_7427929112_200ohm 1 2
Rp 1 2 7190
Cp 1 2 12.644p
Rs 1 N3 0.025
L1 N3 2 8.752u
.ends 1280_7427929112_200ohm
*******
.subckt 1280_7427929115_185ohm 1 2
Rp 1 2 7470
Cp 1 2 9.515p
Rs 1 N3 0.03
L1 N3 2 11.815u
.ends 1280_7427929115_185ohm
*******
